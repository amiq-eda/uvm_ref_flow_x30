/*-------------------------------------------------------------------------
File1 name   : test_lib1.sv
Title1       : Library1 of tests
Project1     :
Created1     :
Description1 : Library1 of tests for the APB1-UART1 Environment1
Notes1       : Includes1 all the test files. Whenever1 a new test case file is 
            : created the file has to be included1 here1
----------------------------------------------------------------------*/
//   Copyright1 1999-2010 Cadence1 Design1 Systems1, Inc1.
//   All Rights1 Reserved1 Worldwide1
//
//   Licensed1 under the Apache1 License1, Version1 2.0 (the
//   "License1"); you may not use this file except1 in
//   compliance1 with the License1.  You may obtain1 a copy of
//   the License1 at
//
//       http1://www1.apache1.org1/licenses1/LICENSE1-2.0
//
//   Unless1 required1 by applicable1 law1 or agreed1 to in
//   writing, software1 distributed1 under the License1 is
//   distributed1 on an "AS1 IS1" BASIS1, WITHOUT1 WARRANTIES1 OR1
//   CONDITIONS1 OF1 ANY1 KIND1, either1 express1 or implied1.  See
//   the License1 for the specific1 language1 governing1
//   permissions1 and limitations1 under the License1.
//----------------------------------------------------------------------

`include "apb_uart_simple_test1.sv"
`include "apb_spi_simple_test1.sv"
`include "apb_gpio_simple_test1.sv"
`include "apb_subsystem_test1.sv"
`include "apb_subsystem_lp_test1.sv"
`include "lp_shutdown_urt11.sv"
