/*-------------------------------------------------------------------------
File19 name   : test_lib19.sv
Title19       : Library19 of tests
Project19     :
Created19     :
Description19 : Library19 of tests for the APB19-UART19 Environment19
Notes19       : Includes19 all the test files. Whenever19 a new test case file is 
            : created the file has to be included19 here19
----------------------------------------------------------------------*/
//   Copyright19 1999-2010 Cadence19 Design19 Systems19, Inc19.
//   All Rights19 Reserved19 Worldwide19
//
//   Licensed19 under the Apache19 License19, Version19 2.0 (the
//   "License19"); you may not use this file except19 in
//   compliance19 with the License19.  You may obtain19 a copy of
//   the License19 at
//
//       http19://www19.apache19.org19/licenses19/LICENSE19-2.0
//
//   Unless19 required19 by applicable19 law19 or agreed19 to in
//   writing, software19 distributed19 under the License19 is
//   distributed19 on an "AS19 IS19" BASIS19, WITHOUT19 WARRANTIES19 OR19
//   CONDITIONS19 OF19 ANY19 KIND19, either19 express19 or implied19.  See
//   the License19 for the specific19 language19 governing19
//   permissions19 and limitations19 under the License19.
//----------------------------------------------------------------------

`include "apb_uart_simple_test19.sv"
`include "apb_spi_simple_test19.sv"
`include "apb_gpio_simple_test19.sv"
`include "apb_subsystem_test19.sv"
`include "apb_subsystem_lp_test19.sv"
`include "lp_shutdown_urt119.sv"
