/*-------------------------------------------------------------------------
File14 name   : uart_internal_if14.sv
Title14       : Interface14 File14
Project14     : UART14 Block Level14
Created14     :
Description14 : Interface14 for collecting14 white14 box14 coverage14
Notes14       :
----------------------------------------------------------------------
Copyright14 2007 (c) Cadence14 Design14 Systems14, Inc14. All Rights14 Reserved14.
----------------------------------------------------------------------*/

interface uart_ctrl_internal_if14(input clock14);
 
  int tx_fifo_ptr14 ;
  int rx_fifo_ptr14 ;

endinterface  
