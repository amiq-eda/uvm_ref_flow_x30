/*-------------------------------------------------------------------------
File9 name   : test_lib9.sv
Title9       : Library9 of tests
Project9     :
Created9     :
Description9 : Library9 of tests for the APB9-UART9 Environment9
Notes9       : Includes9 all the test files. Whenever9 a new test case file is 
            : created the file has to be included9 here9
----------------------------------------------------------------------*/
//   Copyright9 1999-2010 Cadence9 Design9 Systems9, Inc9.
//   All Rights9 Reserved9 Worldwide9
//
//   Licensed9 under the Apache9 License9, Version9 2.0 (the
//   "License9"); you may not use this file except9 in
//   compliance9 with the License9.  You may obtain9 a copy of
//   the License9 at
//
//       http9://www9.apache9.org9/licenses9/LICENSE9-2.0
//
//   Unless9 required9 by applicable9 law9 or agreed9 to in
//   writing, software9 distributed9 under the License9 is
//   distributed9 on an "AS9 IS9" BASIS9, WITHOUT9 WARRANTIES9 OR9
//   CONDITIONS9 OF9 ANY9 KIND9, either9 express9 or implied9.  See
//   the License9 for the specific9 language9 governing9
//   permissions9 and limitations9 under the License9.
//----------------------------------------------------------------------

`include "apb_uart_simple_test9.sv"
`include "apb_spi_simple_test9.sv"
`include "apb_gpio_simple_test9.sv"
`include "apb_subsystem_test9.sv"
`include "apb_subsystem_lp_test9.sv"
`include "lp_shutdown_urt19.sv"
