/*-------------------------------------------------------------------------
File8 name   : test_lib8.sv
Title8       : Library8 of tests
Project8     :
Created8     :
Description8 : Library8 of tests for the APB8-UART8 Environment8
Notes8       : Includes8 all the test files. Whenever8 a new test case file is 
            : created the file has to be included8 here8
----------------------------------------------------------------------*/
//   Copyright8 1999-2010 Cadence8 Design8 Systems8, Inc8.
//   All Rights8 Reserved8 Worldwide8
//
//   Licensed8 under the Apache8 License8, Version8 2.0 (the
//   "License8"); you may not use this file except8 in
//   compliance8 with the License8.  You may obtain8 a copy of
//   the License8 at
//
//       http8://www8.apache8.org8/licenses8/LICENSE8-2.0
//
//   Unless8 required8 by applicable8 law8 or agreed8 to in
//   writing, software8 distributed8 under the License8 is
//   distributed8 on an "AS8 IS8" BASIS8, WITHOUT8 WARRANTIES8 OR8
//   CONDITIONS8 OF8 ANY8 KIND8, either8 express8 or implied8.  See
//   the License8 for the specific8 language8 governing8
//   permissions8 and limitations8 under the License8.
//----------------------------------------------------------------------

`include "apb_uart_simple_test8.sv"
`include "apb_spi_simple_test8.sv"
`include "apb_gpio_simple_test8.sv"
`include "apb_subsystem_test8.sv"
`include "apb_subsystem_lp_test8.sv"
`include "lp_shutdown_urt18.sv"
