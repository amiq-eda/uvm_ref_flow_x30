/*-------------------------------------------------------------------------
File18 name   : test_lib18.sv
Title18       : Library18 of tests
Project18     :
Created18     :
Description18 : Library18 of tests for the APB18-UART18 Environment18
Notes18       : Includes18 all the test files. Whenever18 a new test case file is 
            : created the file has to be included18 here18
----------------------------------------------------------------------*/
//   Copyright18 1999-2010 Cadence18 Design18 Systems18, Inc18.
//   All Rights18 Reserved18 Worldwide18
//
//   Licensed18 under the Apache18 License18, Version18 2.0 (the
//   "License18"); you may not use this file except18 in
//   compliance18 with the License18.  You may obtain18 a copy of
//   the License18 at
//
//       http18://www18.apache18.org18/licenses18/LICENSE18-2.0
//
//   Unless18 required18 by applicable18 law18 or agreed18 to in
//   writing, software18 distributed18 under the License18 is
//   distributed18 on an "AS18 IS18" BASIS18, WITHOUT18 WARRANTIES18 OR18
//   CONDITIONS18 OF18 ANY18 KIND18, either18 express18 or implied18.  See
//   the License18 for the specific18 language18 governing18
//   permissions18 and limitations18 under the License18.
//----------------------------------------------------------------------

`include "apb_uart_simple_test18.sv"
`include "apb_spi_simple_test18.sv"
`include "apb_gpio_simple_test18.sv"
`include "apb_subsystem_test18.sv"
`include "apb_subsystem_lp_test18.sv"
`include "lp_shutdown_urt118.sv"
