/*-------------------------------------------------------------------------
File22 name   : test_lib22.sv
Title22       : Library22 of tests
Project22     :
Created22     :
Description22 : Library22 of tests for the APB22-UART22 Environment22
Notes22       : Includes22 all the test files. Whenever22 a new test case file is 
            : created the file has to be included22 here22
----------------------------------------------------------------------*/
//   Copyright22 1999-2010 Cadence22 Design22 Systems22, Inc22.
//   All Rights22 Reserved22 Worldwide22
//
//   Licensed22 under the Apache22 License22, Version22 2.0 (the
//   "License22"); you may not use this file except22 in
//   compliance22 with the License22.  You may obtain22 a copy of
//   the License22 at
//
//       http22://www22.apache22.org22/licenses22/LICENSE22-2.0
//
//   Unless22 required22 by applicable22 law22 or agreed22 to in
//   writing, software22 distributed22 under the License22 is
//   distributed22 on an "AS22 IS22" BASIS22, WITHOUT22 WARRANTIES22 OR22
//   CONDITIONS22 OF22 ANY22 KIND22, either22 express22 or implied22.  See
//   the License22 for the specific22 language22 governing22
//   permissions22 and limitations22 under the License22.
//----------------------------------------------------------------------

`include "apb_uart_simple_test22.sv"
`include "apb_spi_simple_test22.sv"
`include "apb_gpio_simple_test22.sv"
`include "apb_subsystem_test22.sv"
`include "apb_subsystem_lp_test22.sv"
`include "lp_shutdown_urt122.sv"
