`ifndef AHB_DEFINES23
    `define AHB_DEFINES23

    `ifndef AHB_DATA_WIDTH23
        `define AHB_DATA_WIDTH23 32 // AHB23 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH23
        `define AHB_ADDR_WIDTH23 32 // AHB23 address bus max width
    `endif
`endif
