/*-------------------------------------------------------------------------
File11 name   : spi_defines11.svh
Title11       : APB11 - SPI11 defines11
Project11     :
Created11     :
Description11 : defines11 for the APB11-SPI11 Environment11
Notes11       : 
----------------------------------------------------------------------*/
//   Copyright11 1999-2010 Cadence11 Design11 Systems11, Inc11.
//   All Rights11 Reserved11 Worldwide11
//
//   Licensed11 under the Apache11 License11, Version11 2.0 (the
//   "License11"); you may not use this file except11 in
//   compliance11 with the License11.  You may obtain11 a copy of
//   the License11 at
//
//       http11://www11.apache11.org11/licenses11/LICENSE11-2.0
//
//   Unless11 required11 by applicable11 law11 or agreed11 to in
//   writing, software11 distributed11 under the License11 is
//   distributed11 on an "AS11 IS11" BASIS11, WITHOUT11 WARRANTIES11 OR11
//   CONDITIONS11 OF11 ANY11 KIND11, either11 express11 or implied11.  See
//   the License11 for the specific11 language11 governing11
//   permissions11 and limitations11 under the License11.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH11
`define APB_SPI_DEFINES_SVH11

`define SPI_RX0_REG11    32'h00
`define SPI_RX1_REG11    32'h04
`define SPI_RX2_REG11    32'h08
`define SPI_RX3_REG11    32'h0C
`define SPI_TX0_REG11    32'h00
`define SPI_TX1_REG11    32'h04
`define SPI_TX2_REG11    32'h08
`define SPI_TX3_REG11    32'h0C
`define SPI_CTRL_REG11   32'h10
`define SPI_DIV_REG11    32'h14
`define SPI_SS_REG11     32'h18

`endif
