/*-------------------------------------------------------------------------
File2 name   : spi_defines2.svh
Title2       : APB2 - SPI2 defines2
Project2     :
Created2     :
Description2 : defines2 for the APB2-SPI2 Environment2
Notes2       : 
----------------------------------------------------------------------*/
//   Copyright2 1999-2010 Cadence2 Design2 Systems2, Inc2.
//   All Rights2 Reserved2 Worldwide2
//
//   Licensed2 under the Apache2 License2, Version2 2.0 (the
//   "License2"); you may not use this file except2 in
//   compliance2 with the License2.  You may obtain2 a copy of
//   the License2 at
//
//       http2://www2.apache2.org2/licenses2/LICENSE2-2.0
//
//   Unless2 required2 by applicable2 law2 or agreed2 to in
//   writing, software2 distributed2 under the License2 is
//   distributed2 on an "AS2 IS2" BASIS2, WITHOUT2 WARRANTIES2 OR2
//   CONDITIONS2 OF2 ANY2 KIND2, either2 express2 or implied2.  See
//   the License2 for the specific2 language2 governing2
//   permissions2 and limitations2 under the License2.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH2
`define APB_SPI_DEFINES_SVH2

`define SPI_RX0_REG2    32'h00
`define SPI_RX1_REG2    32'h04
`define SPI_RX2_REG2    32'h08
`define SPI_RX3_REG2    32'h0C
`define SPI_TX0_REG2    32'h00
`define SPI_TX1_REG2    32'h04
`define SPI_TX2_REG2    32'h08
`define SPI_TX3_REG2    32'h0C
`define SPI_CTRL_REG2   32'h10
`define SPI_DIV_REG2    32'h14
`define SPI_SS_REG2     32'h18

`endif
