/*-------------------------------------------------------------------------
File1 name   : spi_defines1.svh
Title1       : APB1 - SPI1 defines1
Project1     :
Created1     :
Description1 : defines1 for the APB1-SPI1 Environment1
Notes1       : 
----------------------------------------------------------------------*/
//   Copyright1 1999-2010 Cadence1 Design1 Systems1, Inc1.
//   All Rights1 Reserved1 Worldwide1
//
//   Licensed1 under the Apache1 License1, Version1 2.0 (the
//   "License1"); you may not use this file except1 in
//   compliance1 with the License1.  You may obtain1 a copy of
//   the License1 at
//
//       http1://www1.apache1.org1/licenses1/LICENSE1-2.0
//
//   Unless1 required1 by applicable1 law1 or agreed1 to in
//   writing, software1 distributed1 under the License1 is
//   distributed1 on an "AS1 IS1" BASIS1, WITHOUT1 WARRANTIES1 OR1
//   CONDITIONS1 OF1 ANY1 KIND1, either1 express1 or implied1.  See
//   the License1 for the specific1 language1 governing1
//   permissions1 and limitations1 under the License1.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH1
`define APB_SPI_DEFINES_SVH1

`define SPI_RX0_REG1    32'h00
`define SPI_RX1_REG1    32'h04
`define SPI_RX2_REG1    32'h08
`define SPI_RX3_REG1    32'h0C
`define SPI_TX0_REG1    32'h00
`define SPI_TX1_REG1    32'h04
`define SPI_TX2_REG1    32'h08
`define SPI_TX3_REG1    32'h0C
`define SPI_CTRL_REG1   32'h10
`define SPI_DIV_REG1    32'h14
`define SPI_SS_REG1     32'h18

`endif
