// IVB23 checksum23: 720351203
/*-----------------------------------------------------------------
File23 name     : ahb_pkg23.sv
Created23       : Wed23 May23 19 15:42:21 2010
Description23   : This23 file imports23 all the files of the OVC23.
Notes23         :
-----------------------------------------------------------------*/
//   Copyright23 1999-2010 Cadence23 Design23 Systems23, Inc23.
//   All Rights23 Reserved23 Worldwide23
//
//   Licensed23 under the Apache23 License23, Version23 2.0 (the
//   "License23"); you may not use this file except23 in
//   compliance23 with the License23.  You may obtain23 a copy of
//   the License23 at
//
//       http23://www23.apache23.org23/licenses23/LICENSE23-2.0
//
//   Unless23 required23 by applicable23 law23 or agreed23 to in
//   writing, software23 distributed23 under the License23 is
//   distributed23 on an "AS23 IS23" BASIS23, WITHOUT23 WARRANTIES23 OR23
//   CONDITIONS23 OF23 ANY23 KIND23, either23 express23 or implied23.  See
//   the License23 for the specific23 language23 governing23
//   permissions23 and limitations23 under the License23.
//----------------------------------------------------------------------


`ifndef AHB_PKG_SV23
`define AHB_PKG_SV23

package ahb_pkg23;

// UVM class library compiled23 in a package
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "ahb_defines23.sv"
`include "ahb_transfer23.sv"

`include "ahb_master_monitor23.sv"
`include "ahb_master_sequencer23.sv"
`include "ahb_master_driver23.sv"
`include "ahb_master_agent23.sv"
// Can23 include universally23 reusable23 master23 sequences here23.

`include "ahb_slave_monitor23.sv"
`include "ahb_slave_sequencer23.sv"
`include "ahb_slave_driver23.sv"
`include "ahb_slave_agent23.sv"
// Can23 include universally23 reusable23 slave23 sequences here23.

`include "ahb_env23.sv"
`include "reg_to_ahb_adapter23.sv"

endpackage : ahb_pkg23

`endif // AHB_PKG_SV23
