/*-------------------------------------------------------------------------
File7 name   : test_lib7.sv
Title7       : Library7 of tests
Project7     :
Created7     :
Description7 : Library7 of tests for the APB7-UART7 Environment7
Notes7       : Includes7 all the test files. Whenever7 a new test case file is 
            : created the file has to be included7 here7
----------------------------------------------------------------------*/
//   Copyright7 1999-2010 Cadence7 Design7 Systems7, Inc7.
//   All Rights7 Reserved7 Worldwide7
//
//   Licensed7 under the Apache7 License7, Version7 2.0 (the
//   "License7"); you may not use this file except7 in
//   compliance7 with the License7.  You may obtain7 a copy of
//   the License7 at
//
//       http7://www7.apache7.org7/licenses7/LICENSE7-2.0
//
//   Unless7 required7 by applicable7 law7 or agreed7 to in
//   writing, software7 distributed7 under the License7 is
//   distributed7 on an "AS7 IS7" BASIS7, WITHOUT7 WARRANTIES7 OR7
//   CONDITIONS7 OF7 ANY7 KIND7, either7 express7 or implied7.  See
//   the License7 for the specific7 language7 governing7
//   permissions7 and limitations7 under the License7.
//----------------------------------------------------------------------

`include "apb_uart_simple_test7.sv"
`include "apb_spi_simple_test7.sv"
`include "apb_gpio_simple_test7.sv"
`include "apb_subsystem_test7.sv"
`include "apb_subsystem_lp_test7.sv"
`include "lp_shutdown_urt17.sv"
