/*-------------------------------------------------------------------------
File13 name   : test_lib13.sv
Title13       : Library13 of tests
Project13     :
Created13     :
Description13 : Library13 of tests for the APB13-UART13 Environment13
Notes13       : Includes13 all the test files. Whenever13 a new test case file is 
            : created the file has to be included13 here13
----------------------------------------------------------------------*/
//   Copyright13 1999-2010 Cadence13 Design13 Systems13, Inc13.
//   All Rights13 Reserved13 Worldwide13
//
//   Licensed13 under the Apache13 License13, Version13 2.0 (the
//   "License13"); you may not use this file except13 in
//   compliance13 with the License13.  You may obtain13 a copy of
//   the License13 at
//
//       http13://www13.apache13.org13/licenses13/LICENSE13-2.0
//
//   Unless13 required13 by applicable13 law13 or agreed13 to in
//   writing, software13 distributed13 under the License13 is
//   distributed13 on an "AS13 IS13" BASIS13, WITHOUT13 WARRANTIES13 OR13
//   CONDITIONS13 OF13 ANY13 KIND13, either13 express13 or implied13.  See
//   the License13 for the specific13 language13 governing13
//   permissions13 and limitations13 under the License13.
//----------------------------------------------------------------------

`include "apb_uart_simple_test13.sv"
`include "apb_spi_simple_test13.sv"
`include "apb_gpio_simple_test13.sv"
`include "apb_subsystem_test13.sv"
`include "apb_subsystem_lp_test13.sv"
`include "lp_shutdown_urt113.sv"
