/*-------------------------------------------------------------------------
File30 name   : spi_defines30.svh
Title30       : APB30 - SPI30 defines30
Project30     :
Created30     :
Description30 : defines30 for the APB30-SPI30 Environment30
Notes30       : 
----------------------------------------------------------------------*/
//   Copyright30 1999-2010 Cadence30 Design30 Systems30, Inc30.
//   All Rights30 Reserved30 Worldwide30
//
//   Licensed30 under the Apache30 License30, Version30 2.0 (the
//   "License30"); you may not use this file except30 in
//   compliance30 with the License30.  You may obtain30 a copy of
//   the License30 at
//
//       http30://www30.apache30.org30/licenses30/LICENSE30-2.0
//
//   Unless30 required30 by applicable30 law30 or agreed30 to in
//   writing, software30 distributed30 under the License30 is
//   distributed30 on an "AS30 IS30" BASIS30, WITHOUT30 WARRANTIES30 OR30
//   CONDITIONS30 OF30 ANY30 KIND30, either30 express30 or implied30.  See
//   the License30 for the specific30 language30 governing30
//   permissions30 and limitations30 under the License30.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH30
`define APB_SPI_DEFINES_SVH30

`define SPI_RX0_REG30    32'h00
`define SPI_RX1_REG30    32'h04
`define SPI_RX2_REG30    32'h08
`define SPI_RX3_REG30    32'h0C
`define SPI_TX0_REG30    32'h00
`define SPI_TX1_REG30    32'h04
`define SPI_TX2_REG30    32'h08
`define SPI_TX3_REG30    32'h0C
`define SPI_CTRL_REG30   32'h10
`define SPI_DIV_REG30    32'h14
`define SPI_SS_REG30     32'h18

`endif
