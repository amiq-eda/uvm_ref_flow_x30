`ifndef AHB_DEFINES28
    `define AHB_DEFINES28

    `ifndef AHB_DATA_WIDTH28
        `define AHB_DATA_WIDTH28 32 // AHB28 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH28
        `define AHB_ADDR_WIDTH28 32 // AHB28 address bus max width
    `endif
`endif
