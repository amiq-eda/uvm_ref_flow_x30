/*-------------------------------------------------------------------------
File27 name   : test_lib27.sv
Title27       : Library27 of tests
Project27     :
Created27     :
Description27 : Library27 of tests for the APB27-UART27 Environment27
Notes27       : Includes27 all the test files. Whenever27 a new test case file is 
            : created the file has to be included27 here27
----------------------------------------------------------------------*/
//   Copyright27 1999-2010 Cadence27 Design27 Systems27, Inc27.
//   All Rights27 Reserved27 Worldwide27
//
//   Licensed27 under the Apache27 License27, Version27 2.0 (the
//   "License27"); you may not use this file except27 in
//   compliance27 with the License27.  You may obtain27 a copy of
//   the License27 at
//
//       http27://www27.apache27.org27/licenses27/LICENSE27-2.0
//
//   Unless27 required27 by applicable27 law27 or agreed27 to in
//   writing, software27 distributed27 under the License27 is
//   distributed27 on an "AS27 IS27" BASIS27, WITHOUT27 WARRANTIES27 OR27
//   CONDITIONS27 OF27 ANY27 KIND27, either27 express27 or implied27.  See
//   the License27 for the specific27 language27 governing27
//   permissions27 and limitations27 under the License27.
//----------------------------------------------------------------------

`include "apb_uart_simple_test27.sv"
`include "apb_spi_simple_test27.sv"
`include "apb_gpio_simple_test27.sv"
`include "apb_subsystem_test27.sv"
`include "apb_subsystem_lp_test27.sv"
`include "lp_shutdown_urt127.sv"
