`ifndef AHB_DEFINES9
    `define AHB_DEFINES9

    `ifndef AHB_DATA_WIDTH9
        `define AHB_DATA_WIDTH9 32 // AHB9 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH9
        `define AHB_ADDR_WIDTH9 32 // AHB9 address bus max width
    `endif
`endif
