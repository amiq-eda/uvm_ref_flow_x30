/*-------------------------------------------------------------------------
File17 name   : gpio_defines17.svh
Title17       : APB17 - GPIO17 defines17
Project17     :
Created17     :
Description17 : defines17 for the APB17-GPIO17 Environment17
Notes17       : 
----------------------------------------------------------------------*/
//   Copyright17 1999-2010 Cadence17 Design17 Systems17, Inc17.
//   All Rights17 Reserved17 Worldwide17
//
//   Licensed17 under the Apache17 License17, Version17 2.0 (the
//   "License17"); you may not use this file except17 in
//   compliance17 with the License17.  You may obtain17 a copy of
//   the License17 at
//
//       http17://www17.apache17.org17/licenses17/LICENSE17-2.0
//
//   Unless17 required17 by applicable17 law17 or agreed17 to in
//   writing, software17 distributed17 under the License17 is
//   distributed17 on an "AS17 IS17" BASIS17, WITHOUT17 WARRANTIES17 OR17
//   CONDITIONS17 OF17 ANY17 KIND17, either17 express17 or implied17.  See
//   the License17 for the specific17 language17 governing17
//   permissions17 and limitations17 under the License17.
//----------------------------------------------------------------------

`ifndef APB_GPIO_DEFINES_SVH17
`define APB_GPIO_DEFINES_SVH17

`define GPIO_DATA_WIDTH17         32
`define GPIO_BYPASS_MODE_REG17    32'h00
`define GPIO_DIRECTION_MODE_REG17 32'h04
`define GPIO_OUTPUT_ENABLE_REG17  32'h08
`define GPIO_OUTPUT_VALUE_REG17   32'h0C
`define GPIO_INPUT_VALUE_REG17    32'h10
`define GPIO_INT_MASK_REG17       32'h14
`define GPIO_INT_ENABLE_REG17     32'h18
`define GPIO_INT_DISABLE_REG17    32'h1C
`define GPIO_INT_STATUS_REG17     32'h20
`define GPIO_INT_TYPE_REG17       32'h24
`define GPIO_INT_VALUE_REG17      32'h28
`define GPIO_INT_ON_ANY_REG17     32'h2C

`endif
