/*-------------------------------------------------------------------------
File4 name   : spi_config4.sv
Title4       : SPI4 environment4 configuration file
Project4     : UVM SystemVerilog4 Cluster4 Level4 Verification4
Created4     :
Description4 :
Notes4       :  
----------------------------------------------------------------------*/
//   Copyright4 1999-2010 Cadence4 Design4 Systems4, Inc4.
//   All Rights4 Reserved4 Worldwide4
//
//   Licensed4 under the Apache4 License4, Version4 2.0 (the
//   "License4"); you may not use this file except4 in
//   compliance4 with the License4.  You may obtain4 a copy of
//   the License4 at
//
//       http4://www4.apache4.org4/licenses4/LICENSE4-2.0
//
//   Unless4 required4 by applicable4 law4 or agreed4 to in
//   writing, software4 distributed4 under the License4 is
//   distributed4 on an "AS4 IS4" BASIS4, WITHOUT4 WARRANTIES4 OR4
//   CONDITIONS4 OF4 ANY4 KIND4, either4 express4 or implied4.  See
//   the License4 for the specific4 language4 governing4
//   permissions4 and limitations4 under the License4.
//----------------------------------------------------------------------


`ifndef SPI_CFG_SVH4
`define SPI_CFG_SVH4

class spi_config4 extends uvm_object;

  function new (string name = "");
    super.new(name);
  endfunction

  uvm_active_passive_enum  active_passive4 = UVM_ACTIVE;

  `uvm_object_utils_begin(spi_config4)
    `uvm_field_enum(uvm_active_passive_enum, active_passive4, UVM_ALL_ON)
   `uvm_object_utils_end

endclass

`endif

