`ifndef AHB_DEFINES6
    `define AHB_DEFINES6

    `ifndef AHB_DATA_WIDTH6
        `define AHB_DATA_WIDTH6 32 // AHB6 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH6
        `define AHB_ADDR_WIDTH6 32 // AHB6 address bus max width
    `endif
`endif
