// IVB15 checksum15: 720351203
/*-----------------------------------------------------------------
File15 name     : ahb_pkg15.sv
Created15       : Wed15 May15 19 15:42:21 2010
Description15   : This15 file imports15 all the files of the OVC15.
Notes15         :
-----------------------------------------------------------------*/
//   Copyright15 1999-2010 Cadence15 Design15 Systems15, Inc15.
//   All Rights15 Reserved15 Worldwide15
//
//   Licensed15 under the Apache15 License15, Version15 2.0 (the
//   "License15"); you may not use this file except15 in
//   compliance15 with the License15.  You may obtain15 a copy of
//   the License15 at
//
//       http15://www15.apache15.org15/licenses15/LICENSE15-2.0
//
//   Unless15 required15 by applicable15 law15 or agreed15 to in
//   writing, software15 distributed15 under the License15 is
//   distributed15 on an "AS15 IS15" BASIS15, WITHOUT15 WARRANTIES15 OR15
//   CONDITIONS15 OF15 ANY15 KIND15, either15 express15 or implied15.  See
//   the License15 for the specific15 language15 governing15
//   permissions15 and limitations15 under the License15.
//----------------------------------------------------------------------


`ifndef AHB_PKG_SV15
`define AHB_PKG_SV15

package ahb_pkg15;

// UVM class library compiled15 in a package
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "ahb_defines15.sv"
`include "ahb_transfer15.sv"

`include "ahb_master_monitor15.sv"
`include "ahb_master_sequencer15.sv"
`include "ahb_master_driver15.sv"
`include "ahb_master_agent15.sv"
// Can15 include universally15 reusable15 master15 sequences here15.

`include "ahb_slave_monitor15.sv"
`include "ahb_slave_sequencer15.sv"
`include "ahb_slave_driver15.sv"
`include "ahb_slave_agent15.sv"
// Can15 include universally15 reusable15 slave15 sequences here15.

`include "ahb_env15.sv"
`include "reg_to_ahb_adapter15.sv"

endpackage : ahb_pkg15

`endif // AHB_PKG_SV15
