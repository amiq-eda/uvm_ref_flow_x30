`ifndef AHB_DEFINES24
    `define AHB_DEFINES24

    `ifndef AHB_DATA_WIDTH24
        `define AHB_DATA_WIDTH24 32 // AHB24 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH24
        `define AHB_ADDR_WIDTH24 32 // AHB24 address bus max width
    `endif
`endif
