/*-------------------------------------------------------------------------
File2 name   : test_lib2.sv
Title2       : Library2 of tests
Project2     :
Created2     :
Description2 : Library2 of tests for the APB2-UART2 Environment2
Notes2       : Includes2 all the test files. Whenever2 a new test case file is 
            : created the file has to be included2 here2
----------------------------------------------------------------------*/
//   Copyright2 1999-2010 Cadence2 Design2 Systems2, Inc2.
//   All Rights2 Reserved2 Worldwide2
//
//   Licensed2 under the Apache2 License2, Version2 2.0 (the
//   "License2"); you may not use this file except2 in
//   compliance2 with the License2.  You may obtain2 a copy of
//   the License2 at
//
//       http2://www2.apache2.org2/licenses2/LICENSE2-2.0
//
//   Unless2 required2 by applicable2 law2 or agreed2 to in
//   writing, software2 distributed2 under the License2 is
//   distributed2 on an "AS2 IS2" BASIS2, WITHOUT2 WARRANTIES2 OR2
//   CONDITIONS2 OF2 ANY2 KIND2, either2 express2 or implied2.  See
//   the License2 for the specific2 language2 governing2
//   permissions2 and limitations2 under the License2.
//----------------------------------------------------------------------

`include "apb_uart_simple_test2.sv"
`include "apb_spi_simple_test2.sv"
`include "apb_gpio_simple_test2.sv"
`include "apb_subsystem_test2.sv"
`include "apb_subsystem_lp_test2.sv"
`include "lp_shutdown_urt12.sv"
