/*-------------------------------------------------------------------------
File1 name   : uart_ctrl_virtual_sequencer1.sv
Title1       : Virtual sequencer
Project1     :
Created1     :
Description1 : This1 file implements1 the Virtual sequencer for APB1-UART1 environment1
Notes1       : 
----------------------------------------------------------------------*/
//   Copyright1 1999-2010 Cadence1 Design1 Systems1, Inc1.
//   All Rights1 Reserved1 Worldwide1
//
//   Licensed1 under the Apache1 License1, Version1 2.0 (the
//   "License1"); you may not use this file except1 in
//   compliance1 with the License1.  You may obtain1 a copy of
//   the License1 at
//
//       http1://www1.apache1.org1/licenses1/LICENSE1-2.0
//
//   Unless1 required1 by applicable1 law1 or agreed1 to in
//   writing, software1 distributed1 under the License1 is
//   distributed1 on an "AS1 IS1" BASIS1, WITHOUT1 WARRANTIES1 OR1
//   CONDITIONS1 OF1 ANY1 KIND1, either1 express1 or implied1.  See
//   the License1 for the specific1 language1 governing1
//   permissions1 and limitations1 under the License1.
//----------------------------------------------------------------------


class uart_ctrl_virtual_sequencer1 extends uvm_sequencer;

    apb_pkg1::apb_master_sequencer1 apb_seqr1;
    uart_pkg1::uart_sequencer1 uart_seqr1;
    uart_ctrl_reg_sequencer1 reg_seqr;

    // UVM_REG: Pointer1 to the register model
    uart_ctrl_reg_model_c1 reg_model1;
   
    // Uart1 Controller1 configuration object
    uart_ctrl_config1 cfg;

    function new (input string name="uart_ctrl_virtual_sequencer1", input uvm_component parent=null);
      super.new(name, parent);
    endfunction : new

    `uvm_component_utils_begin(uart_ctrl_virtual_sequencer1)
       `uvm_field_object(cfg, UVM_DEFAULT | UVM_NOPRINT)
       `uvm_field_object(reg_model1, UVM_DEFAULT | UVM_REFERENCE)
    `uvm_component_utils_end

endclass : uart_ctrl_virtual_sequencer1
