`ifndef AHB_DEFINES4
    `define AHB_DEFINES4

    `ifndef AHB_DATA_WIDTH4
        `define AHB_DATA_WIDTH4 32 // AHB4 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH4
        `define AHB_ADDR_WIDTH4 32 // AHB4 address bus max width
    `endif
`endif
