/*-------------------------------------------------------------------------
File17 name   : spi_defines17.svh
Title17       : APB17 - SPI17 defines17
Project17     :
Created17     :
Description17 : defines17 for the APB17-SPI17 Environment17
Notes17       : 
----------------------------------------------------------------------*/
//   Copyright17 1999-2010 Cadence17 Design17 Systems17, Inc17.
//   All Rights17 Reserved17 Worldwide17
//
//   Licensed17 under the Apache17 License17, Version17 2.0 (the
//   "License17"); you may not use this file except17 in
//   compliance17 with the License17.  You may obtain17 a copy of
//   the License17 at
//
//       http17://www17.apache17.org17/licenses17/LICENSE17-2.0
//
//   Unless17 required17 by applicable17 law17 or agreed17 to in
//   writing, software17 distributed17 under the License17 is
//   distributed17 on an "AS17 IS17" BASIS17, WITHOUT17 WARRANTIES17 OR17
//   CONDITIONS17 OF17 ANY17 KIND17, either17 express17 or implied17.  See
//   the License17 for the specific17 language17 governing17
//   permissions17 and limitations17 under the License17.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH17
`define APB_SPI_DEFINES_SVH17

`define SPI_RX0_REG17    32'h00
`define SPI_RX1_REG17    32'h04
`define SPI_RX2_REG17    32'h08
`define SPI_RX3_REG17    32'h0C
`define SPI_TX0_REG17    32'h00
`define SPI_TX1_REG17    32'h04
`define SPI_TX2_REG17    32'h08
`define SPI_TX3_REG17    32'h0C
`define SPI_CTRL_REG17   32'h10
`define SPI_DIV_REG17    32'h14
`define SPI_SS_REG17     32'h18

`endif
