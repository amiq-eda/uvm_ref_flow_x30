`ifndef AHB_DEFINES3
    `define AHB_DEFINES3

    `ifndef AHB_DATA_WIDTH3
        `define AHB_DATA_WIDTH3 32 // AHB3 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH3
        `define AHB_ADDR_WIDTH3 32 // AHB3 address bus max width
    `endif
`endif
