`ifndef AHB_DEFINES8
    `define AHB_DEFINES8

    `ifndef AHB_DATA_WIDTH8
        `define AHB_DATA_WIDTH8 32 // AHB8 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH8
        `define AHB_ADDR_WIDTH8 32 // AHB8 address bus max width
    `endif
`endif
