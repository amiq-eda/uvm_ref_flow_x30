`ifndef AHB_DEFINES1
    `define AHB_DEFINES1

    `ifndef AHB_DATA_WIDTH1
        `define AHB_DATA_WIDTH1 32 // AHB1 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH1
        `define AHB_ADDR_WIDTH1 32 // AHB1 address bus max width
    `endif
`endif
