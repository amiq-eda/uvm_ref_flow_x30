/*-------------------------------------------------------------------------
File30 name   : test_lib30.sv
Title30       : Library30 of tests
Project30     :
Created30     :
Description30 : Library30 of tests for the APB30-UART30 Environment30
Notes30       : Includes30 all the test files. Whenever30 a new test case file is 
            : created the file has to be included30 here30
----------------------------------------------------------------------*/
//   Copyright30 1999-2010 Cadence30 Design30 Systems30, Inc30.
//   All Rights30 Reserved30 Worldwide30
//
//   Licensed30 under the Apache30 License30, Version30 2.0 (the
//   "License30"); you may not use this file except30 in
//   compliance30 with the License30.  You may obtain30 a copy of
//   the License30 at
//
//       http30://www30.apache30.org30/licenses30/LICENSE30-2.0
//
//   Unless30 required30 by applicable30 law30 or agreed30 to in
//   writing, software30 distributed30 under the License30 is
//   distributed30 on an "AS30 IS30" BASIS30, WITHOUT30 WARRANTIES30 OR30
//   CONDITIONS30 OF30 ANY30 KIND30, either30 express30 or implied30.  See
//   the License30 for the specific30 language30 governing30
//   permissions30 and limitations30 under the License30.
//----------------------------------------------------------------------

`include "apb_uart_simple_test30.sv"
`include "apb_spi_simple_test30.sv"
`include "apb_gpio_simple_test30.sv"
`include "apb_subsystem_test30.sv"
`include "apb_subsystem_lp_test30.sv"
`include "lp_shutdown_urt130.sv"
