/*-------------------------------------------------------------------------
File28 name   : uart_internal_if28.sv
Title28       : Interface28 File28
Project28     : UART28 Block Level28
Created28     :
Description28 : Interface28 for collecting28 white28 box28 coverage28
Notes28       :
----------------------------------------------------------------------
Copyright28 2007 (c) Cadence28 Design28 Systems28, Inc28. All Rights28 Reserved28.
----------------------------------------------------------------------*/

interface uart_ctrl_internal_if28(input clock28);
 
  int tx_fifo_ptr28 ;
  int rx_fifo_ptr28 ;

endinterface  
