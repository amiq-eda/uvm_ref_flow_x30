`ifndef AHB_DEFINES5
    `define AHB_DEFINES5

    `ifndef AHB_DATA_WIDTH5
        `define AHB_DATA_WIDTH5 32 // AHB5 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH5
        `define AHB_ADDR_WIDTH5 32 // AHB5 address bus max width
    `endif
`endif
