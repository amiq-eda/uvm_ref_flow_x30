`ifndef AHB_DEFINES17
    `define AHB_DEFINES17

    `ifndef AHB_DATA_WIDTH17
        `define AHB_DATA_WIDTH17 32 // AHB17 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH17
        `define AHB_ADDR_WIDTH17 32 // AHB17 address bus max width
    `endif
`endif
