/*-------------------------------------------------------------------------
File23 name   : test_lib23.sv
Title23       : Library23 of tests
Project23     :
Created23     :
Description23 : Library23 of tests for the APB23-UART23 Environment23
Notes23       : Includes23 all the test files. Whenever23 a new test case file is 
            : created the file has to be included23 here23
----------------------------------------------------------------------*/
//   Copyright23 1999-2010 Cadence23 Design23 Systems23, Inc23.
//   All Rights23 Reserved23 Worldwide23
//
//   Licensed23 under the Apache23 License23, Version23 2.0 (the
//   "License23"); you may not use this file except23 in
//   compliance23 with the License23.  You may obtain23 a copy of
//   the License23 at
//
//       http23://www23.apache23.org23/licenses23/LICENSE23-2.0
//
//   Unless23 required23 by applicable23 law23 or agreed23 to in
//   writing, software23 distributed23 under the License23 is
//   distributed23 on an "AS23 IS23" BASIS23, WITHOUT23 WARRANTIES23 OR23
//   CONDITIONS23 OF23 ANY23 KIND23, either23 express23 or implied23.  See
//   the License23 for the specific23 language23 governing23
//   permissions23 and limitations23 under the License23.
//----------------------------------------------------------------------

`include "apb_uart_simple_test23.sv"
`include "apb_spi_simple_test23.sv"
`include "apb_gpio_simple_test23.sv"
`include "apb_subsystem_test23.sv"
`include "apb_subsystem_lp_test23.sv"
`include "lp_shutdown_urt123.sv"
