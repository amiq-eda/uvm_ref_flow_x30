/*-------------------------------------------------------------------------
File4 name   : test_lib4.sv
Title4       : Library4 of tests
Project4     :
Created4     :
Description4 : Library4 of tests for the APB4-UART4 Environment4
Notes4       : Includes4 all the test files. Whenever4 a new test case file is 
            : created the file has to be included4 here4
----------------------------------------------------------------------*/
//   Copyright4 1999-2010 Cadence4 Design4 Systems4, Inc4.
//   All Rights4 Reserved4 Worldwide4
//
//   Licensed4 under the Apache4 License4, Version4 2.0 (the
//   "License4"); you may not use this file except4 in
//   compliance4 with the License4.  You may obtain4 a copy of
//   the License4 at
//
//       http4://www4.apache4.org4/licenses4/LICENSE4-2.0
//
//   Unless4 required4 by applicable4 law4 or agreed4 to in
//   writing, software4 distributed4 under the License4 is
//   distributed4 on an "AS4 IS4" BASIS4, WITHOUT4 WARRANTIES4 OR4
//   CONDITIONS4 OF4 ANY4 KIND4, either4 express4 or implied4.  See
//   the License4 for the specific4 language4 governing4
//   permissions4 and limitations4 under the License4.
//----------------------------------------------------------------------

`include "apb_uart_simple_test4.sv"
`include "apb_spi_simple_test4.sv"
`include "apb_gpio_simple_test4.sv"
`include "apb_subsystem_test4.sv"
`include "apb_subsystem_lp_test4.sv"
`include "lp_shutdown_urt14.sv"
