/*-------------------------------------------------------------------------
File7 name   : spi_defines7.svh
Title7       : APB7 - SPI7 defines7
Project7     :
Created7     :
Description7 : defines7 for the APB7-SPI7 Environment7
Notes7       : 
----------------------------------------------------------------------*/
//   Copyright7 1999-2010 Cadence7 Design7 Systems7, Inc7.
//   All Rights7 Reserved7 Worldwide7
//
//   Licensed7 under the Apache7 License7, Version7 2.0 (the
//   "License7"); you may not use this file except7 in
//   compliance7 with the License7.  You may obtain7 a copy of
//   the License7 at
//
//       http7://www7.apache7.org7/licenses7/LICENSE7-2.0
//
//   Unless7 required7 by applicable7 law7 or agreed7 to in
//   writing, software7 distributed7 under the License7 is
//   distributed7 on an "AS7 IS7" BASIS7, WITHOUT7 WARRANTIES7 OR7
//   CONDITIONS7 OF7 ANY7 KIND7, either7 express7 or implied7.  See
//   the License7 for the specific7 language7 governing7
//   permissions7 and limitations7 under the License7.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH7
`define APB_SPI_DEFINES_SVH7

`define SPI_RX0_REG7    32'h00
`define SPI_RX1_REG7    32'h04
`define SPI_RX2_REG7    32'h08
`define SPI_RX3_REG7    32'h0C
`define SPI_TX0_REG7    32'h00
`define SPI_TX1_REG7    32'h04
`define SPI_TX2_REG7    32'h08
`define SPI_TX3_REG7    32'h0C
`define SPI_CTRL_REG7   32'h10
`define SPI_DIV_REG7    32'h14
`define SPI_SS_REG7     32'h18

`endif
