/*-------------------------------------------------------------------------
File17 name   : test_lib17.sv
Title17       : Library17 of tests
Project17     :
Created17     :
Description17 : Library17 of tests for the APB17-UART17 Environment17
Notes17       : Includes17 all the test files. Whenever17 a new test case file is 
            : created the file has to be included17 here17
----------------------------------------------------------------------*/
//   Copyright17 1999-2010 Cadence17 Design17 Systems17, Inc17.
//   All Rights17 Reserved17 Worldwide17
//
//   Licensed17 under the Apache17 License17, Version17 2.0 (the
//   "License17"); you may not use this file except17 in
//   compliance17 with the License17.  You may obtain17 a copy of
//   the License17 at
//
//       http17://www17.apache17.org17/licenses17/LICENSE17-2.0
//
//   Unless17 required17 by applicable17 law17 or agreed17 to in
//   writing, software17 distributed17 under the License17 is
//   distributed17 on an "AS17 IS17" BASIS17, WITHOUT17 WARRANTIES17 OR17
//   CONDITIONS17 OF17 ANY17 KIND17, either17 express17 or implied17.  See
//   the License17 for the specific17 language17 governing17
//   permissions17 and limitations17 under the License17.
//----------------------------------------------------------------------

`include "apb_uart_simple_test17.sv"
`include "apb_spi_simple_test17.sv"
`include "apb_gpio_simple_test17.sv"
`include "apb_subsystem_test17.sv"
`include "apb_subsystem_lp_test17.sv"
`include "lp_shutdown_urt117.sv"
