`ifndef AHB_DEFINES30
    `define AHB_DEFINES30

    `ifndef AHB_DATA_WIDTH30
        `define AHB_DATA_WIDTH30 32 // AHB30 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH30
        `define AHB_ADDR_WIDTH30 32 // AHB30 address bus max width
    `endif
`endif
