/*-------------------------------------------------------------------------
File11 name   : test_lib11.sv
Title11       : Library11 of tests
Project11     :
Created11     :
Description11 : Library11 of tests for the APB11-UART11 Environment11
Notes11       : Includes11 all the test files. Whenever11 a new test case file is 
            : created the file has to be included11 here11
----------------------------------------------------------------------*/
//   Copyright11 1999-2010 Cadence11 Design11 Systems11, Inc11.
//   All Rights11 Reserved11 Worldwide11
//
//   Licensed11 under the Apache11 License11, Version11 2.0 (the
//   "License11"); you may not use this file except11 in
//   compliance11 with the License11.  You may obtain11 a copy of
//   the License11 at
//
//       http11://www11.apache11.org11/licenses11/LICENSE11-2.0
//
//   Unless11 required11 by applicable11 law11 or agreed11 to in
//   writing, software11 distributed11 under the License11 is
//   distributed11 on an "AS11 IS11" BASIS11, WITHOUT11 WARRANTIES11 OR11
//   CONDITIONS11 OF11 ANY11 KIND11, either11 express11 or implied11.  See
//   the License11 for the specific11 language11 governing11
//   permissions11 and limitations11 under the License11.
//----------------------------------------------------------------------

`include "apb_uart_simple_test11.sv"
`include "apb_spi_simple_test11.sv"
`include "apb_gpio_simple_test11.sv"
`include "apb_subsystem_test11.sv"
`include "apb_subsystem_lp_test11.sv"
`include "lp_shutdown_urt111.sv"
