/*-------------------------------------------------------------------------
File27 name   : spi_defines27.svh
Title27       : APB27 - SPI27 defines27
Project27     :
Created27     :
Description27 : defines27 for the APB27-SPI27 Environment27
Notes27       : 
----------------------------------------------------------------------*/
//   Copyright27 1999-2010 Cadence27 Design27 Systems27, Inc27.
//   All Rights27 Reserved27 Worldwide27
//
//   Licensed27 under the Apache27 License27, Version27 2.0 (the
//   "License27"); you may not use this file except27 in
//   compliance27 with the License27.  You may obtain27 a copy of
//   the License27 at
//
//       http27://www27.apache27.org27/licenses27/LICENSE27-2.0
//
//   Unless27 required27 by applicable27 law27 or agreed27 to in
//   writing, software27 distributed27 under the License27 is
//   distributed27 on an "AS27 IS27" BASIS27, WITHOUT27 WARRANTIES27 OR27
//   CONDITIONS27 OF27 ANY27 KIND27, either27 express27 or implied27.  See
//   the License27 for the specific27 language27 governing27
//   permissions27 and limitations27 under the License27.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH27
`define APB_SPI_DEFINES_SVH27

`define SPI_RX0_REG27    32'h00
`define SPI_RX1_REG27    32'h04
`define SPI_RX2_REG27    32'h08
`define SPI_RX3_REG27    32'h0C
`define SPI_TX0_REG27    32'h00
`define SPI_TX1_REG27    32'h04
`define SPI_TX2_REG27    32'h08
`define SPI_TX3_REG27    32'h0C
`define SPI_CTRL_REG27   32'h10
`define SPI_DIV_REG27    32'h14
`define SPI_SS_REG27     32'h18

`endif
