`ifndef AHB_DEFINES16
    `define AHB_DEFINES16

    `ifndef AHB_DATA_WIDTH16
        `define AHB_DATA_WIDTH16 32 // AHB16 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH16
        `define AHB_ADDR_WIDTH16 32 // AHB16 address bus max width
    `endif
`endif
