/*-------------------------------------------------------------------------
File14 name   : spi_defines14.svh
Title14       : APB14 - SPI14 defines14
Project14     :
Created14     :
Description14 : defines14 for the APB14-SPI14 Environment14
Notes14       : 
----------------------------------------------------------------------*/
//   Copyright14 1999-2010 Cadence14 Design14 Systems14, Inc14.
//   All Rights14 Reserved14 Worldwide14
//
//   Licensed14 under the Apache14 License14, Version14 2.0 (the
//   "License14"); you may not use this file except14 in
//   compliance14 with the License14.  You may obtain14 a copy of
//   the License14 at
//
//       http14://www14.apache14.org14/licenses14/LICENSE14-2.0
//
//   Unless14 required14 by applicable14 law14 or agreed14 to in
//   writing, software14 distributed14 under the License14 is
//   distributed14 on an "AS14 IS14" BASIS14, WITHOUT14 WARRANTIES14 OR14
//   CONDITIONS14 OF14 ANY14 KIND14, either14 express14 or implied14.  See
//   the License14 for the specific14 language14 governing14
//   permissions14 and limitations14 under the License14.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH14
`define APB_SPI_DEFINES_SVH14

`define SPI_RX0_REG14    32'h00
`define SPI_RX1_REG14    32'h04
`define SPI_RX2_REG14    32'h08
`define SPI_RX3_REG14    32'h0C
`define SPI_TX0_REG14    32'h00
`define SPI_TX1_REG14    32'h04
`define SPI_TX2_REG14    32'h08
`define SPI_TX3_REG14    32'h0C
`define SPI_CTRL_REG14   32'h10
`define SPI_DIV_REG14    32'h14
`define SPI_SS_REG14     32'h18

`endif
