/*-------------------------------------------------------------------------
File10 name   : test_lib10.sv
Title10       : Library10 of tests
Project10     :
Created10     :
Description10 : Library10 of tests for the APB10-UART10 Environment10
Notes10       : Includes10 all the test files. Whenever10 a new test case file is 
            : created the file has to be included10 here10
----------------------------------------------------------------------*/
//   Copyright10 1999-2010 Cadence10 Design10 Systems10, Inc10.
//   All Rights10 Reserved10 Worldwide10
//
//   Licensed10 under the Apache10 License10, Version10 2.0 (the
//   "License10"); you may not use this file except10 in
//   compliance10 with the License10.  You may obtain10 a copy of
//   the License10 at
//
//       http10://www10.apache10.org10/licenses10/LICENSE10-2.0
//
//   Unless10 required10 by applicable10 law10 or agreed10 to in
//   writing, software10 distributed10 under the License10 is
//   distributed10 on an "AS10 IS10" BASIS10, WITHOUT10 WARRANTIES10 OR10
//   CONDITIONS10 OF10 ANY10 KIND10, either10 express10 or implied10.  See
//   the License10 for the specific10 language10 governing10
//   permissions10 and limitations10 under the License10.
//----------------------------------------------------------------------

`include "apb_uart_simple_test10.sv"
`include "apb_spi_simple_test10.sv"
`include "apb_gpio_simple_test10.sv"
`include "apb_subsystem_test10.sv"
`include "apb_subsystem_lp_test10.sv"
`include "lp_shutdown_urt110.sv"
