`ifndef AHB_DEFINES22
    `define AHB_DEFINES22

    `ifndef AHB_DATA_WIDTH22
        `define AHB_DATA_WIDTH22 32 // AHB22 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH22
        `define AHB_ADDR_WIDTH22 32 // AHB22 address bus max width
    `endif
`endif
