/*-------------------------------------------------------------------------
File26 name   : test_lib26.sv
Title26       : Library26 of tests
Project26     :
Created26     :
Description26 : Library26 of tests for the APB26-UART26 Environment26
Notes26       : Includes26 all the test files. Whenever26 a new test case file is 
            : created the file has to be included26 here26
----------------------------------------------------------------------*/
//   Copyright26 1999-2010 Cadence26 Design26 Systems26, Inc26.
//   All Rights26 Reserved26 Worldwide26
//
//   Licensed26 under the Apache26 License26, Version26 2.0 (the
//   "License26"); you may not use this file except26 in
//   compliance26 with the License26.  You may obtain26 a copy of
//   the License26 at
//
//       http26://www26.apache26.org26/licenses26/LICENSE26-2.0
//
//   Unless26 required26 by applicable26 law26 or agreed26 to in
//   writing, software26 distributed26 under the License26 is
//   distributed26 on an "AS26 IS26" BASIS26, WITHOUT26 WARRANTIES26 OR26
//   CONDITIONS26 OF26 ANY26 KIND26, either26 express26 or implied26.  See
//   the License26 for the specific26 language26 governing26
//   permissions26 and limitations26 under the License26.
//----------------------------------------------------------------------

`include "apb_uart_simple_test26.sv"
`include "apb_spi_simple_test26.sv"
`include "apb_gpio_simple_test26.sv"
`include "apb_subsystem_test26.sv"
`include "apb_subsystem_lp_test26.sv"
`include "lp_shutdown_urt126.sv"
