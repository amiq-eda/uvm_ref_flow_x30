/*-------------------------------------------------------------------------
File24 name   : test_lib24.sv
Title24       : Library24 of tests
Project24     :
Created24     :
Description24 : Library24 of tests for the APB24-UART24 Environment24
Notes24       : Includes24 all the test files. Whenever24 a new test case file is 
            : created the file has to be included24 here24
----------------------------------------------------------------------*/
//   Copyright24 1999-2010 Cadence24 Design24 Systems24, Inc24.
//   All Rights24 Reserved24 Worldwide24
//
//   Licensed24 under the Apache24 License24, Version24 2.0 (the
//   "License24"); you may not use this file except24 in
//   compliance24 with the License24.  You may obtain24 a copy of
//   the License24 at
//
//       http24://www24.apache24.org24/licenses24/LICENSE24-2.0
//
//   Unless24 required24 by applicable24 law24 or agreed24 to in
//   writing, software24 distributed24 under the License24 is
//   distributed24 on an "AS24 IS24" BASIS24, WITHOUT24 WARRANTIES24 OR24
//   CONDITIONS24 OF24 ANY24 KIND24, either24 express24 or implied24.  See
//   the License24 for the specific24 language24 governing24
//   permissions24 and limitations24 under the License24.
//----------------------------------------------------------------------

`include "apb_uart_simple_test24.sv"
`include "apb_spi_simple_test24.sv"
`include "apb_gpio_simple_test24.sv"
`include "apb_subsystem_test24.sv"
`include "apb_subsystem_lp_test24.sv"
`include "lp_shutdown_urt124.sv"
