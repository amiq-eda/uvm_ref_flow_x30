/*-------------------------------------------------------------------------
File29 name   : uart_internal_if29.sv
Title29       : Interface29 File29
Project29     : UART29 Block Level29
Created29     :
Description29 : Interface29 for collecting29 white29 box29 coverage29
Notes29       :
----------------------------------------------------------------------
Copyright29 2007 (c) Cadence29 Design29 Systems29, Inc29. All Rights29 Reserved29.
----------------------------------------------------------------------*/

interface uart_ctrl_internal_if29(input clock29);
 
  int tx_fifo_ptr29 ;
  int rx_fifo_ptr29 ;

endinterface  
