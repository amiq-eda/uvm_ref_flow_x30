`ifndef AHB_DEFINES2
    `define AHB_DEFINES2

    `ifndef AHB_DATA_WIDTH2
        `define AHB_DATA_WIDTH2 32 // AHB2 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH2
        `define AHB_ADDR_WIDTH2 32 // AHB2 address bus max width
    `endif
`endif
