/*-------------------------------------------------------------------------
File17 name   : uart_internal_if17.sv
Title17       : Interface17 File17
Project17     : UART17 Block Level17
Created17     :
Description17 : Interface17 for collecting17 white17 box17 coverage17
Notes17       :
----------------------------------------------------------------------
Copyright17 2007 (c) Cadence17 Design17 Systems17, Inc17. All Rights17 Reserved17.
----------------------------------------------------------------------*/

interface uart_ctrl_internal_if17(input clock17);
 
  int tx_fifo_ptr17 ;
  int rx_fifo_ptr17 ;

endinterface  
