`ifndef AHB_DEFINES15
    `define AHB_DEFINES15

    `ifndef AHB_DATA_WIDTH15
        `define AHB_DATA_WIDTH15 32 // AHB15 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH15
        `define AHB_ADDR_WIDTH15 32 // AHB15 address bus max width
    `endif
`endif
