/*-------------------------------------------------------------------------
File9 name   : gpio_if9.sv
Title9       : GPIO9 SystemVerilog9 UVM UVC9
Project9     : SystemVerilog9 UVM Cluster9 Level9 Verification9
Created9     :
Description9 : 
Notes9       :  
---------------------------------------------------------------------------*/
//   Copyright9 1999-2010 Cadence9 Design9 Systems9, Inc9.
//   All Rights9 Reserved9 Worldwide9
//
//   Licensed9 under the Apache9 License9, Version9 2.0 (the
//   "License9"); you may not use this file except9 in
//   compliance9 with the License9.  You may obtain9 a copy of
//   the License9 at
//
//       http9://www9.apache9.org9/licenses9/LICENSE9-2.0
//
//   Unless9 required9 by applicable9 law9 or agreed9 to in
//   writing, software9 distributed9 under the License9 is
//   distributed9 on an "AS9 IS9" BASIS9, WITHOUT9 WARRANTIES9 OR9
//   CONDITIONS9 OF9 ANY9 KIND9, either9 express9 or implied9.  See
//   the License9 for the specific9 language9 governing9
//   permissions9 and limitations9 under the License9.
//----------------------------------------------------------------------


interface gpio_if9();

  // Control9 flags9
  bit                has_checks9 = 1;
  bit                has_coverage = 1;

  // Actual9 Signals9
  // APB9 Slave9 Interface9 - inputs9
  logic              pclk9;
  logic              n_p_reset9;

  // Slave9 GPIO9 Interface9 - inputs9
  logic [`GPIO_DATA_WIDTH9-1:0]       n_gpio_pin_oe9;
  logic [`GPIO_DATA_WIDTH9-1:0]       gpio_pin_out9;
  logic [`GPIO_DATA_WIDTH9-1:0]       gpio_pin_in9;

// Coverage9 and assertions9 to be implemented here9.

/*
always @(negedge sig_pclk9)
begin

// Read and write never true9 at the same time
assertReadOrWrite9: assert property (
                   disable iff(!has_checks9) 
                   ($onehot(sig_grant9) |-> !(sig_read9 && sig_write9)))
                   else
                     $error("ERR_READ_OR_WRITE9\n Read and Write true9 at \
                             the same time");

end
*/

endinterface : gpio_if9

