/*-------------------------------------------------------------------------
File25 name   : test_lib25.sv
Title25       : Library25 of tests
Project25     :
Created25     :
Description25 : Library25 of tests for the APB25-UART25 Environment25
Notes25       : Includes25 all the test files. Whenever25 a new test case file is 
            : created the file has to be included25 here25
----------------------------------------------------------------------*/
//   Copyright25 1999-2010 Cadence25 Design25 Systems25, Inc25.
//   All Rights25 Reserved25 Worldwide25
//
//   Licensed25 under the Apache25 License25, Version25 2.0 (the
//   "License25"); you may not use this file except25 in
//   compliance25 with the License25.  You may obtain25 a copy of
//   the License25 at
//
//       http25://www25.apache25.org25/licenses25/LICENSE25-2.0
//
//   Unless25 required25 by applicable25 law25 or agreed25 to in
//   writing, software25 distributed25 under the License25 is
//   distributed25 on an "AS25 IS25" BASIS25, WITHOUT25 WARRANTIES25 OR25
//   CONDITIONS25 OF25 ANY25 KIND25, either25 express25 or implied25.  See
//   the License25 for the specific25 language25 governing25
//   permissions25 and limitations25 under the License25.
//----------------------------------------------------------------------

`include "apb_uart_simple_test25.sv"
`include "apb_spi_simple_test25.sv"
`include "apb_gpio_simple_test25.sv"
`include "apb_subsystem_test25.sv"
`include "apb_subsystem_lp_test25.sv"
`include "lp_shutdown_urt125.sv"
