`ifndef SPI_RDB_SV16
`define SPI_RDB_SV16

// Input16 File16: spi_rgm16.spirit16

// Number16 of addrMaps16 = 1
// Number16 of regFiles16 = 1
// Number16 of registers = 3
// Number16 of memories = 0


//////////////////////////////////////////////////////////////////////////////
// Register definition16
//////////////////////////////////////////////////////////////////////////////
// Line16 Number16: 23


class spi_ctrl_c16 extends uvm_reg;

  rand uvm_reg_field char_len16;
  rand uvm_reg_field go_bsy16;
  rand uvm_reg_field rx_neg16;
  rand uvm_reg_field tx_neg16;
  rand uvm_reg_field lsb;
  rand uvm_reg_field ie16;
  rand uvm_reg_field ass16;

  constraint c_char_len16 { char_len16.value == 7'b0001000; }
  constraint c_tx_neg16 { tx_neg16.value == 1'b1; }
  constraint c_rx_neg16 { rx_neg16.value == 1'b1; }
  constraint c_lsb16 { lsb.value == 1'b1; }
  constraint c_ie16 { ie16.value == 1'b1; }
  constraint c_ass16 { ass16.value == 1'b1; }
  virtual function void build();
    char_len16 = uvm_reg_field::type_id::create("char_len16");
    char_len16.configure(this, 7, 0, "RW", 0, `UVM_REG_DATA_WIDTH'h0>>0, 1, 1, 1);
    go_bsy16 = uvm_reg_field::type_id::create("go_bsy16");
    go_bsy16.configure(this, 1, 8, "RW", 0, `UVM_REG_DATA_WIDTH'h0>>8, 1, 1, 1);
    rx_neg16 = uvm_reg_field::type_id::create("rx_neg16");
    rx_neg16.configure(this, 1, 9, "RW", 0, `UVM_REG_DATA_WIDTH'h0>>9, 1, 1, 1);
    tx_neg16 = uvm_reg_field::type_id::create("tx_neg16");
    tx_neg16.configure(this, 1, 10, "RW", 0, `UVM_REG_DATA_WIDTH'h0>>10, 1, 1, 1);
    lsb = uvm_reg_field::type_id::create("lsb");
    lsb.configure(this, 1, 11, "RW", 0, `UVM_REG_DATA_WIDTH'h0>>11, 1, 1, 1);
    ie16 = uvm_reg_field::type_id::create("ie16");
    ie16.configure(this, 1, 12, "RW", 0, `UVM_REG_DATA_WIDTH'h0>>12, 1, 1, 1);
    ass16 = uvm_reg_field::type_id::create("ass16");
    ass16.configure(this, 1, 13, "RW", 0, `UVM_REG_DATA_WIDTH'h0>>13, 1, 1, 1);
  endfunction

  covergroup value_cg16;
    option.per_instance=1;
    coverpoint char_len16.value[6:0];
    coverpoint go_bsy16.value[0:0];
    coverpoint rx_neg16.value[0:0];
    coverpoint tx_neg16.value[0:0];
    coverpoint lsb.value[0:0];
    coverpoint ie16.value[0:0];
    coverpoint ass16.value[0:0];
  endgroup
  
  virtual function void sample_values();
    super.sample_values();
    value_cg16.sample();
  endfunction

  `uvm_register_cb(spi_ctrl_c16, uvm_reg_cbs) 
  `uvm_set_super_type(spi_ctrl_c16, uvm_reg)
  `uvm_object_utils(spi_ctrl_c16)
  function new(input string name="unnamed16-spi_ctrl_c16");
    super.new(name, 32, build_coverage(UVM_CVR_FIELD_VALS));
    if(has_coverage(UVM_CVR_FIELD_VALS)) value_cg16=new;
  endfunction : new
endclass : spi_ctrl_c16

//////////////////////////////////////////////////////////////////////////////
// Register definition16
//////////////////////////////////////////////////////////////////////////////
// Line16 Number16: 99


class spi_divider_c16 extends uvm_reg;

  rand uvm_reg_field divider16;

  constraint c_divider16 { divider16.value == 16'b1; }
  virtual function void build();
    divider16 = uvm_reg_field::type_id::create("divider16");
    divider16.configure(this, 16, 0, "RW", 0, `UVM_REG_DATA_WIDTH'hffff>>0, 1, 1, 1);
  endfunction

  covergroup value_cg16;
    option.per_instance=1;
    coverpoint divider16.value[15:0];
  endgroup
  
  virtual function void sample_values();
    super.sample_values();
    value_cg16.sample();
  endfunction

  `uvm_register_cb(spi_divider_c16, uvm_reg_cbs) 
  `uvm_set_super_type(spi_divider_c16, uvm_reg)
  `uvm_object_utils(spi_divider_c16)
  function new(input string name="unnamed16-spi_divider_c16");
    super.new(name, 32, build_coverage(UVM_CVR_FIELD_VALS));
    if(has_coverage(UVM_CVR_FIELD_VALS)) value_cg16=new;
  endfunction : new
endclass : spi_divider_c16

//////////////////////////////////////////////////////////////////////////////
// Register definition16
//////////////////////////////////////////////////////////////////////////////
// Line16 Number16: 122


class spi_ss_c16 extends uvm_reg;

  rand uvm_reg_field ss;

  constraint c_ss16 { ss.value == 8'b1; }
  virtual function void build();
    ss = uvm_reg_field::type_id::create("ss");
    ss.configure(this, 8, 0, "RW", 0, `UVM_REG_DATA_WIDTH'h0>>0, 1, 1, 1);
  endfunction

  covergroup value_cg16;
    option.per_instance=1;
    coverpoint ss.value[7:0];
  endgroup
  
  virtual function void sample_values();
    super.sample_values();
    value_cg16.sample();
  endfunction

  `uvm_register_cb(spi_ss_c16, uvm_reg_cbs) 
  `uvm_set_super_type(spi_ss_c16, uvm_reg)
  `uvm_object_utils(spi_ss_c16)
  function new(input string name="unnamed16-spi_ss_c16");
    super.new(name, 32, build_coverage(UVM_CVR_FIELD_VALS));
    if(has_coverage(UVM_CVR_FIELD_VALS)) value_cg16=new;
  endfunction : new
endclass : spi_ss_c16

class spi_regfile16 extends uvm_reg_block;

  rand spi_ctrl_c16 spi_ctrl16;
  rand spi_divider_c16 spi_divider16;
  rand spi_ss_c16 spi_ss16;

  virtual function void build();

    // Now16 create all registers

    spi_ctrl16 = spi_ctrl_c16::type_id::create("spi_ctrl16", , get_full_name());
    spi_divider16 = spi_divider_c16::type_id::create("spi_divider16", , get_full_name());
    spi_ss16 = spi_ss_c16::type_id::create("spi_ss16", , get_full_name());

    // Now16 build the registers. Set parent and hdl_paths

    spi_ctrl16.configure(this, null, "spi_ctrl_reg16");
    spi_ctrl16.build();
    spi_divider16.configure(this, null, "spi_divider_reg16");
    spi_divider16.build();
    spi_ss16.configure(this, null, "spi_ss_reg16");
    spi_ss16.build();
    // Now16 define address mappings16
    default_map = create_map("default_map", 0, 4, UVM_LITTLE_ENDIAN);
    default_map.add_reg(spi_ctrl16, `UVM_REG_ADDR_WIDTH'h10, "RW");
    default_map.add_reg(spi_divider16, `UVM_REG_ADDR_WIDTH'h14, "RW");
    default_map.add_reg(spi_ss16, `UVM_REG_ADDR_WIDTH'h18, "RW");
  endfunction

  `uvm_object_utils(spi_regfile16)
  function new(input string name="unnamed16-spi_rf16");
    super.new(name, UVM_NO_COVERAGE);
  endfunction : new
endclass : spi_regfile16

//////////////////////////////////////////////////////////////////////////////
// Address_map16 definition16
//////////////////////////////////////////////////////////////////////////////
class spi_reg_model_c16 extends uvm_reg_block;

  rand spi_regfile16 spi_rf16;

  function void build();
    // Now16 define address mappings16
    default_map = create_map("default_map", 0, 4, UVM_LITTLE_ENDIAN);
    spi_rf16 = spi_regfile16::type_id::create("spi_rf16", , get_full_name());
    spi_rf16.configure(this, "rf216");
    spi_rf16.build();
    spi_rf16.lock_model();
    default_map.add_submap(spi_rf16.default_map, `UVM_REG_ADDR_WIDTH'h800000);
    set_hdl_path_root("apb_spi_addr_map_c16");
    this.lock_model();
  endfunction
  `uvm_object_utils(spi_reg_model_c16)
  function new(input string name="unnamed16-spi_reg_model_c16");
    super.new(name, UVM_NO_COVERAGE);
  endfunction
endclass : spi_reg_model_c16

`endif // SPI_RDB_SV16
