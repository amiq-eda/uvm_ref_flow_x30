/*-------------------------------------------------------------------------
File24 name   : spi_defines24.svh
Title24       : APB24 - SPI24 defines24
Project24     :
Created24     :
Description24 : defines24 for the APB24-SPI24 Environment24
Notes24       : 
----------------------------------------------------------------------*/
//   Copyright24 1999-2010 Cadence24 Design24 Systems24, Inc24.
//   All Rights24 Reserved24 Worldwide24
//
//   Licensed24 under the Apache24 License24, Version24 2.0 (the
//   "License24"); you may not use this file except24 in
//   compliance24 with the License24.  You may obtain24 a copy of
//   the License24 at
//
//       http24://www24.apache24.org24/licenses24/LICENSE24-2.0
//
//   Unless24 required24 by applicable24 law24 or agreed24 to in
//   writing, software24 distributed24 under the License24 is
//   distributed24 on an "AS24 IS24" BASIS24, WITHOUT24 WARRANTIES24 OR24
//   CONDITIONS24 OF24 ANY24 KIND24, either24 express24 or implied24.  See
//   the License24 for the specific24 language24 governing24
//   permissions24 and limitations24 under the License24.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH24
`define APB_SPI_DEFINES_SVH24

`define SPI_RX0_REG24    32'h00
`define SPI_RX1_REG24    32'h04
`define SPI_RX2_REG24    32'h08
`define SPI_RX3_REG24    32'h0C
`define SPI_TX0_REG24    32'h00
`define SPI_TX1_REG24    32'h04
`define SPI_TX2_REG24    32'h08
`define SPI_TX3_REG24    32'h0C
`define SPI_CTRL_REG24   32'h10
`define SPI_DIV_REG24    32'h14
`define SPI_SS_REG24     32'h18

`endif
