/*-------------------------------------------------------------------------
File1 name   : uart_internal_if1.sv
Title1       : Interface1 File1
Project1     : UART1 Block Level1
Created1     :
Description1 : Interface1 for collecting1 white1 box1 coverage1
Notes1       :
----------------------------------------------------------------------
Copyright1 2007 (c) Cadence1 Design1 Systems1, Inc1. All Rights1 Reserved1.
----------------------------------------------------------------------*/

interface uart_ctrl_internal_if1(input clock1);
 
  int tx_fifo_ptr1 ;
  int rx_fifo_ptr1 ;

endinterface  
