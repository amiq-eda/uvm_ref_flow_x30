`ifndef AHB_DEFINES29
    `define AHB_DEFINES29

    `ifndef AHB_DATA_WIDTH29
        `define AHB_DATA_WIDTH29 32 // AHB29 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH29
        `define AHB_ADDR_WIDTH29 32 // AHB29 address bus max width
    `endif
`endif
