/*-------------------------------------------------------------------------
File18 name   : uart_internal_if18.sv
Title18       : Interface18 File18
Project18     : UART18 Block Level18
Created18     :
Description18 : Interface18 for collecting18 white18 box18 coverage18
Notes18       :
----------------------------------------------------------------------
Copyright18 2007 (c) Cadence18 Design18 Systems18, Inc18. All Rights18 Reserved18.
----------------------------------------------------------------------*/

interface uart_ctrl_internal_if18(input clock18);
 
  int tx_fifo_ptr18 ;
  int rx_fifo_ptr18 ;

endinterface  
