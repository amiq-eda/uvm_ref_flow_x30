/*-------------------------------------------------------------------------
File1 name   : apb_subsystem_vir_sequencer1.sv
Title1       : Virtual sequencer
Project1     :
Created1     :
Description1 : This1 file implements1 the Virtual sequencer for APB1-UART1 environment1
Notes1       : 
----------------------------------------------------------------------*/
//   Copyright1 1999-2010 Cadence1 Design1 Systems1, Inc1.
//   All Rights1 Reserved1 Worldwide1
//
//   Licensed1 under the Apache1 License1, Version1 2.0 (the
//   "License1"); you may not use this file except1 in
//   compliance1 with the License1.  You may obtain1 a copy of
//   the License1 at
//
//       http1://www1.apache1.org1/licenses1/LICENSE1-2.0
//
//   Unless1 required1 by applicable1 law1 or agreed1 to in
//   writing, software1 distributed1 under the License1 is
//   distributed1 on an "AS1 IS1" BASIS1, WITHOUT1 WARRANTIES1 OR1
//   CONDITIONS1 OF1 ANY1 KIND1, either1 express1 or implied1.  See
//   the License1 for the specific1 language1 governing1
//   permissions1 and limitations1 under the License1.
//----------------------------------------------------------------------

class apb_subsystem_virtual_sequencer1 extends uvm_sequencer;

    ahb_pkg1::ahb_master_sequencer1 ahb_seqr1;
    uart_pkg1::uart_sequencer1 uart0_seqr1;
    uart_pkg1::uart_sequencer1 uart1_seqr1;
    spi_sequencer1 spi0_seqr1;
    gpio_sequencer1 gpio0_seqr1;
    apb_ss_reg_model_c1 reg_model_ptr1;
    
    function new (string name, uvm_component parent);
      super.new(name, parent);
    endfunction : new

    `uvm_component_utils_begin(apb_subsystem_virtual_sequencer1)
       `uvm_field_object(reg_model_ptr1, UVM_DEFAULT | UVM_REFERENCE)
    `uvm_component_utils_end

endclass : apb_subsystem_virtual_sequencer1

