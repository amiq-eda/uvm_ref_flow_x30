`ifndef AHB_DEFINES25
    `define AHB_DEFINES25

    `ifndef AHB_DATA_WIDTH25
        `define AHB_DATA_WIDTH25 32 // AHB25 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH25
        `define AHB_ADDR_WIDTH25 32 // AHB25 address bus max width
    `endif
`endif
