`ifndef AHB_DEFINES14
    `define AHB_DEFINES14

    `ifndef AHB_DATA_WIDTH14
        `define AHB_DATA_WIDTH14 32 // AHB14 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH14
        `define AHB_ADDR_WIDTH14 32 // AHB14 address bus max width
    `endif
`endif
