/*-------------------------------------------------------------------------
File28 name   : test_lib28.sv
Title28       : Library28 of tests
Project28     :
Created28     :
Description28 : Library28 of tests for the APB28-UART28 Environment28
Notes28       : Includes28 all the test files. Whenever28 a new test case file is 
            : created the file has to be included28 here28
----------------------------------------------------------------------*/
//   Copyright28 1999-2010 Cadence28 Design28 Systems28, Inc28.
//   All Rights28 Reserved28 Worldwide28
//
//   Licensed28 under the Apache28 License28, Version28 2.0 (the
//   "License28"); you may not use this file except28 in
//   compliance28 with the License28.  You may obtain28 a copy of
//   the License28 at
//
//       http28://www28.apache28.org28/licenses28/LICENSE28-2.0
//
//   Unless28 required28 by applicable28 law28 or agreed28 to in
//   writing, software28 distributed28 under the License28 is
//   distributed28 on an "AS28 IS28" BASIS28, WITHOUT28 WARRANTIES28 OR28
//   CONDITIONS28 OF28 ANY28 KIND28, either28 express28 or implied28.  See
//   the License28 for the specific28 language28 governing28
//   permissions28 and limitations28 under the License28.
//----------------------------------------------------------------------

`include "apb_uart_simple_test28.sv"
`include "apb_spi_simple_test28.sv"
`include "apb_gpio_simple_test28.sv"
`include "apb_subsystem_test28.sv"
`include "apb_subsystem_lp_test28.sv"
`include "lp_shutdown_urt128.sv"
