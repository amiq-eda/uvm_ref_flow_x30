/*-------------------------------------------------------------------------
File15 name   : spi_defines15.svh
Title15       : APB15 - SPI15 defines15
Project15     :
Created15     :
Description15 : defines15 for the APB15-SPI15 Environment15
Notes15       : 
----------------------------------------------------------------------*/
//   Copyright15 1999-2010 Cadence15 Design15 Systems15, Inc15.
//   All Rights15 Reserved15 Worldwide15
//
//   Licensed15 under the Apache15 License15, Version15 2.0 (the
//   "License15"); you may not use this file except15 in
//   compliance15 with the License15.  You may obtain15 a copy of
//   the License15 at
//
//       http15://www15.apache15.org15/licenses15/LICENSE15-2.0
//
//   Unless15 required15 by applicable15 law15 or agreed15 to in
//   writing, software15 distributed15 under the License15 is
//   distributed15 on an "AS15 IS15" BASIS15, WITHOUT15 WARRANTIES15 OR15
//   CONDITIONS15 OF15 ANY15 KIND15, either15 express15 or implied15.  See
//   the License15 for the specific15 language15 governing15
//   permissions15 and limitations15 under the License15.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH15
`define APB_SPI_DEFINES_SVH15

`define SPI_RX0_REG15    32'h00
`define SPI_RX1_REG15    32'h04
`define SPI_RX2_REG15    32'h08
`define SPI_RX3_REG15    32'h0C
`define SPI_TX0_REG15    32'h00
`define SPI_TX1_REG15    32'h04
`define SPI_TX2_REG15    32'h08
`define SPI_TX3_REG15    32'h0C
`define SPI_CTRL_REG15   32'h10
`define SPI_DIV_REG15    32'h14
`define SPI_SS_REG15     32'h18

`endif
