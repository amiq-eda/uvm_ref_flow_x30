/*-------------------------------------------------------------------------
File25 name   : spi_defines25.svh
Title25       : APB25 - SPI25 defines25
Project25     :
Created25     :
Description25 : defines25 for the APB25-SPI25 Environment25
Notes25       : 
----------------------------------------------------------------------*/
//   Copyright25 1999-2010 Cadence25 Design25 Systems25, Inc25.
//   All Rights25 Reserved25 Worldwide25
//
//   Licensed25 under the Apache25 License25, Version25 2.0 (the
//   "License25"); you may not use this file except25 in
//   compliance25 with the License25.  You may obtain25 a copy of
//   the License25 at
//
//       http25://www25.apache25.org25/licenses25/LICENSE25-2.0
//
//   Unless25 required25 by applicable25 law25 or agreed25 to in
//   writing, software25 distributed25 under the License25 is
//   distributed25 on an "AS25 IS25" BASIS25, WITHOUT25 WARRANTIES25 OR25
//   CONDITIONS25 OF25 ANY25 KIND25, either25 express25 or implied25.  See
//   the License25 for the specific25 language25 governing25
//   permissions25 and limitations25 under the License25.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH25
`define APB_SPI_DEFINES_SVH25

`define SPI_RX0_REG25    32'h00
`define SPI_RX1_REG25    32'h04
`define SPI_RX2_REG25    32'h08
`define SPI_RX3_REG25    32'h0C
`define SPI_TX0_REG25    32'h00
`define SPI_TX1_REG25    32'h04
`define SPI_TX2_REG25    32'h08
`define SPI_TX3_REG25    32'h0C
`define SPI_CTRL_REG25   32'h10
`define SPI_DIV_REG25    32'h14
`define SPI_SS_REG25     32'h18

`endif
