/*-------------------------------------------------------------------------
File9 name   : spi_defines9.svh
Title9       : APB9 - SPI9 defines9
Project9     :
Created9     :
Description9 : defines9 for the APB9-SPI9 Environment9
Notes9       : 
----------------------------------------------------------------------*/
//   Copyright9 1999-2010 Cadence9 Design9 Systems9, Inc9.
//   All Rights9 Reserved9 Worldwide9
//
//   Licensed9 under the Apache9 License9, Version9 2.0 (the
//   "License9"); you may not use this file except9 in
//   compliance9 with the License9.  You may obtain9 a copy of
//   the License9 at
//
//       http9://www9.apache9.org9/licenses9/LICENSE9-2.0
//
//   Unless9 required9 by applicable9 law9 or agreed9 to in
//   writing, software9 distributed9 under the License9 is
//   distributed9 on an "AS9 IS9" BASIS9, WITHOUT9 WARRANTIES9 OR9
//   CONDITIONS9 OF9 ANY9 KIND9, either9 express9 or implied9.  See
//   the License9 for the specific9 language9 governing9
//   permissions9 and limitations9 under the License9.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH9
`define APB_SPI_DEFINES_SVH9

`define SPI_RX0_REG9    32'h00
`define SPI_RX1_REG9    32'h04
`define SPI_RX2_REG9    32'h08
`define SPI_RX3_REG9    32'h0C
`define SPI_TX0_REG9    32'h00
`define SPI_TX1_REG9    32'h04
`define SPI_TX2_REG9    32'h08
`define SPI_TX3_REG9    32'h0C
`define SPI_CTRL_REG9   32'h10
`define SPI_DIV_REG9    32'h14
`define SPI_SS_REG9     32'h18

`endif
