/*-------------------------------------------------------------------------
File10 name   : apb_pkg10.sv
Title10       : Package10 for APB10 UVC10
Project10     :
Created10     :
Description10 : 
Notes10       :  
----------------------------------------------------------------------*/
//   Copyright10 1999-2010 Cadence10 Design10 Systems10, Inc10.
//   All Rights10 Reserved10 Worldwide10
//
//   Licensed10 under the Apache10 License10, Version10 2.0 (the
//   "License10"); you may not use this file except10 in
//   compliance10 with the License10.  You may obtain10 a copy of
//   the License10 at
//
//       http10://www10.apache10.org10/licenses10/LICENSE10-2.0
//
//   Unless10 required10 by applicable10 law10 or agreed10 to in
//   writing, software10 distributed10 under the License10 is
//   distributed10 on an "AS10 IS10" BASIS10, WITHOUT10 WARRANTIES10 OR10
//   CONDITIONS10 OF10 ANY10 KIND10, either10 express10 or implied10.  See
//   the License10 for the specific10 language10 governing10
//   permissions10 and limitations10 under the License10.
//----------------------------------------------------------------------

  
`ifndef APB_PKG_SV10
`define APB_PKG_SV10

package apb_pkg10;

// Import10 the UVM class library  and UVM automation10 macros10
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "apb_config10.sv"
`include "apb_types10.sv"
`include "apb_transfer10.sv"
`include "apb_monitor10.sv"
`include "apb_collector10.sv"

`include "apb_master_driver10.sv"
`include "apb_master_sequencer10.sv"
`include "apb_master_agent10.sv"

`include "apb_slave_driver10.sv"
`include "apb_slave_sequencer10.sv"
`include "apb_slave_agent10.sv"

`include "apb_master_seq_lib10.sv"
`include "apb_slave_seq_lib10.sv"

`include "apb_env10.sv"

`include "reg_to_apb_adapter10.sv"

endpackage : apb_pkg10
`endif  // APB_PKG_SV10
