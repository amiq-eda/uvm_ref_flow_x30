/*-------------------------------------------------------------------------
File6 name   : test_lib6.sv
Title6       : Library6 of tests
Project6     :
Created6     :
Description6 : Library6 of tests for the APB6-UART6 Environment6
Notes6       : Includes6 all the test files. Whenever6 a new test case file is 
            : created the file has to be included6 here6
----------------------------------------------------------------------*/
//   Copyright6 1999-2010 Cadence6 Design6 Systems6, Inc6.
//   All Rights6 Reserved6 Worldwide6
//
//   Licensed6 under the Apache6 License6, Version6 2.0 (the
//   "License6"); you may not use this file except6 in
//   compliance6 with the License6.  You may obtain6 a copy of
//   the License6 at
//
//       http6://www6.apache6.org6/licenses6/LICENSE6-2.0
//
//   Unless6 required6 by applicable6 law6 or agreed6 to in
//   writing, software6 distributed6 under the License6 is
//   distributed6 on an "AS6 IS6" BASIS6, WITHOUT6 WARRANTIES6 OR6
//   CONDITIONS6 OF6 ANY6 KIND6, either6 express6 or implied6.  See
//   the License6 for the specific6 language6 governing6
//   permissions6 and limitations6 under the License6.
//----------------------------------------------------------------------

`include "apb_uart_simple_test6.sv"
`include "apb_spi_simple_test6.sv"
`include "apb_gpio_simple_test6.sv"
`include "apb_subsystem_test6.sv"
`include "apb_subsystem_lp_test6.sv"
`include "lp_shutdown_urt16.sv"
