/*-------------------------------------------------------------------------
File22 name   : spi_defines22.svh
Title22       : APB22 - SPI22 defines22
Project22     :
Created22     :
Description22 : defines22 for the APB22-SPI22 Environment22
Notes22       : 
----------------------------------------------------------------------*/
//   Copyright22 1999-2010 Cadence22 Design22 Systems22, Inc22.
//   All Rights22 Reserved22 Worldwide22
//
//   Licensed22 under the Apache22 License22, Version22 2.0 (the
//   "License22"); you may not use this file except22 in
//   compliance22 with the License22.  You may obtain22 a copy of
//   the License22 at
//
//       http22://www22.apache22.org22/licenses22/LICENSE22-2.0
//
//   Unless22 required22 by applicable22 law22 or agreed22 to in
//   writing, software22 distributed22 under the License22 is
//   distributed22 on an "AS22 IS22" BASIS22, WITHOUT22 WARRANTIES22 OR22
//   CONDITIONS22 OF22 ANY22 KIND22, either22 express22 or implied22.  See
//   the License22 for the specific22 language22 governing22
//   permissions22 and limitations22 under the License22.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH22
`define APB_SPI_DEFINES_SVH22

`define SPI_RX0_REG22    32'h00
`define SPI_RX1_REG22    32'h04
`define SPI_RX2_REG22    32'h08
`define SPI_RX3_REG22    32'h0C
`define SPI_TX0_REG22    32'h00
`define SPI_TX1_REG22    32'h04
`define SPI_TX2_REG22    32'h08
`define SPI_TX3_REG22    32'h0C
`define SPI_CTRL_REG22   32'h10
`define SPI_DIV_REG22    32'h14
`define SPI_SS_REG22     32'h18

`endif
