/*-------------------------------------------------------------------------
File12 name   : test_lib12.sv
Title12       : Library12 of tests
Project12     :
Created12     :
Description12 : Library12 of tests for the APB12-UART12 Environment12
Notes12       : Includes12 all the test files. Whenever12 a new test case file is 
            : created the file has to be included12 here12
----------------------------------------------------------------------*/
//   Copyright12 1999-2010 Cadence12 Design12 Systems12, Inc12.
//   All Rights12 Reserved12 Worldwide12
//
//   Licensed12 under the Apache12 License12, Version12 2.0 (the
//   "License12"); you may not use this file except12 in
//   compliance12 with the License12.  You may obtain12 a copy of
//   the License12 at
//
//       http12://www12.apache12.org12/licenses12/LICENSE12-2.0
//
//   Unless12 required12 by applicable12 law12 or agreed12 to in
//   writing, software12 distributed12 under the License12 is
//   distributed12 on an "AS12 IS12" BASIS12, WITHOUT12 WARRANTIES12 OR12
//   CONDITIONS12 OF12 ANY12 KIND12, either12 express12 or implied12.  See
//   the License12 for the specific12 language12 governing12
//   permissions12 and limitations12 under the License12.
//----------------------------------------------------------------------

`include "apb_uart_simple_test12.sv"
`include "apb_spi_simple_test12.sv"
`include "apb_gpio_simple_test12.sv"
`include "apb_subsystem_test12.sv"
`include "apb_subsystem_lp_test12.sv"
`include "lp_shutdown_urt112.sv"
