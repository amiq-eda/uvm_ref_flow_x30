/*-------------------------------------------------------------------------
File5 name   : test_lib5.sv
Title5       : Library5 of tests
Project5     :
Created5     :
Description5 : Library5 of tests for the APB5-UART5 Environment5
Notes5       : Includes5 all the test files. Whenever5 a new test case file is 
            : created the file has to be included5 here5
----------------------------------------------------------------------*/
//   Copyright5 1999-2010 Cadence5 Design5 Systems5, Inc5.
//   All Rights5 Reserved5 Worldwide5
//
//   Licensed5 under the Apache5 License5, Version5 2.0 (the
//   "License5"); you may not use this file except5 in
//   compliance5 with the License5.  You may obtain5 a copy of
//   the License5 at
//
//       http5://www5.apache5.org5/licenses5/LICENSE5-2.0
//
//   Unless5 required5 by applicable5 law5 or agreed5 to in
//   writing, software5 distributed5 under the License5 is
//   distributed5 on an "AS5 IS5" BASIS5, WITHOUT5 WARRANTIES5 OR5
//   CONDITIONS5 OF5 ANY5 KIND5, either5 express5 or implied5.  See
//   the License5 for the specific5 language5 governing5
//   permissions5 and limitations5 under the License5.
//----------------------------------------------------------------------

`include "apb_uart_simple_test5.sv"
`include "apb_spi_simple_test5.sv"
`include "apb_gpio_simple_test5.sv"
`include "apb_subsystem_test5.sv"
`include "apb_subsystem_lp_test5.sv"
`include "lp_shutdown_urt15.sv"
