// This14 file is generated14 using Cadence14 iregGen14 version14 1.05

`ifndef UART_CTRL_REGS_SV14
`define UART_CTRL_REGS_SV14

// Input14 File14: uart_ctrl_regs14.xml14

// Number14 of AddrMaps14 = 1
// Number14 of RegFiles14 = 1
// Number14 of Registers14 = 6
// Number14 of Memories14 = 0


//////////////////////////////////////////////////////////////////////////////
// Register definition14
//////////////////////////////////////////////////////////////////////////////
// Line14 Number14: 262


class ua_div_latch0_c14 extends uvm_reg;

  rand uvm_reg_field div_val14;

  constraint c_div_val14 { div_val14.value == 1; }
  virtual function void build();
    div_val14 = uvm_reg_field::type_id::create("div_val14");
    div_val14.configure(this, 8, 0, "RW", 0, `UVM_REG_DATA_WIDTH'h00>>0, 1, 1, 1);
    wr_cg14.set_inst_name($sformatf("%s.wcov14", get_full_name()));
    rd_cg14.set_inst_name($sformatf("%s.rcov14", get_full_name()));
  endfunction

  covergroup wr_cg14;
    option.per_instance=1;
    div_val14 : coverpoint div_val14.value[7:0];
  endgroup
  covergroup rd_cg14;
    option.per_instance=1;
    div_val14 : coverpoint div_val14.value[7:0];
  endgroup

  virtual function void sample(uvm_reg_data_t  data, byte_en, bit is_read, uvm_reg_map map);
    super.sample(data, byte_en, is_read, map);
    if(!is_read) wr_cg14.sample();
    if(is_read) rd_cg14.sample();
  endfunction

  `uvm_register_cb(ua_div_latch0_c14, uvm_reg_cbs) 
  `uvm_set_super_type(ua_div_latch0_c14, uvm_reg)
  `uvm_object_utils(ua_div_latch0_c14)
  function new(input string name="unnamed14-ua_div_latch0_c14");
    super.new(name, 8, build_coverage(UVM_CVR_FIELD_VALS));
    wr_cg14=new;
    rd_cg14=new;
  endfunction : new
endclass : ua_div_latch0_c14

//////////////////////////////////////////////////////////////////////////////
// Register definition14
//////////////////////////////////////////////////////////////////////////////
// Line14 Number14: 287


class ua_div_latch1_c14 extends uvm_reg;

  rand uvm_reg_field div_val14;

  constraint c_div_val14 { div_val14.value == 0; }
  virtual function void build();
    div_val14 = uvm_reg_field::type_id::create("div_val14");
    div_val14.configure(this, 8, 0, "RW", 0, `UVM_REG_DATA_WIDTH'h00>>0, 1, 1, 1);
    wr_cg14.set_inst_name($sformatf("%s.wcov14", get_full_name()));
    rd_cg14.set_inst_name($sformatf("%s.rcov14", get_full_name()));
  endfunction

  covergroup wr_cg14;
    option.per_instance=1;
    div_val14 : coverpoint div_val14.value[7:0];
  endgroup
  covergroup rd_cg14;
    option.per_instance=1;
    div_val14 : coverpoint div_val14.value[7:0];
  endgroup

  virtual function void sample(uvm_reg_data_t  data, byte_en, bit is_read, uvm_reg_map map);
    super.sample(data, byte_en, is_read, map);
    if(!is_read) wr_cg14.sample();
    if(is_read) rd_cg14.sample();
  endfunction

  `uvm_register_cb(ua_div_latch1_c14, uvm_reg_cbs) 
  `uvm_set_super_type(ua_div_latch1_c14, uvm_reg)
  `uvm_object_utils(ua_div_latch1_c14)
  function new(input string name="unnamed14-ua_div_latch1_c14");
    super.new(name, 8, build_coverage(UVM_CVR_FIELD_VALS));
    wr_cg14=new;
    rd_cg14=new;
  endfunction : new
endclass : ua_div_latch1_c14

//////////////////////////////////////////////////////////////////////////////
// Register definition14
//////////////////////////////////////////////////////////////////////////////
// Line14 Number14: 82


class ua_int_id_c14 extends uvm_reg;

  uvm_reg_field priority_bit14;
  uvm_reg_field bit114;
  uvm_reg_field bit214;
  uvm_reg_field bit314;

  virtual function void build();
    priority_bit14 = uvm_reg_field::type_id::create("priority_bit14");
    priority_bit14.configure(this, 1, 0, "RO", 0, `UVM_REG_DATA_WIDTH'hC1>>0, 1, 0, 1);
    bit114 = uvm_reg_field::type_id::create("bit114");
    bit114.configure(this, 1, 1, "RO", 0, `UVM_REG_DATA_WIDTH'hC1>>1, 1, 0, 1);
    bit214 = uvm_reg_field::type_id::create("bit214");
    bit214.configure(this, 1, 2, "RO", 0, `UVM_REG_DATA_WIDTH'hC1>>2, 1, 0, 1);
    bit314 = uvm_reg_field::type_id::create("bit314");
    bit314.configure(this, 1, 3, "RO", 0, `UVM_REG_DATA_WIDTH'hC1>>3, 1, 0, 1);
    rd_cg14.set_inst_name($sformatf("%s.rcov14", get_full_name()));
  endfunction

  covergroup rd_cg14;
    option.per_instance=1;
    priority_bit14 : coverpoint priority_bit14.value[0:0];
    bit114 : coverpoint bit114.value[0:0];
    bit214 : coverpoint bit214.value[0:0];
    bit314 : coverpoint bit314.value[0:0];
  endgroup

  virtual function void sample(uvm_reg_data_t  data, byte_en, bit is_read, uvm_reg_map map);
    super.sample(data, byte_en, is_read, map);
    if(is_read) rd_cg14.sample();
  endfunction

  `uvm_register_cb(ua_int_id_c14, uvm_reg_cbs) 
  `uvm_set_super_type(ua_int_id_c14, uvm_reg)
  `uvm_object_utils(ua_int_id_c14)
  function new(input string name="unnamed14-ua_int_id_c14");
    super.new(name, 8, build_coverage(UVM_CVR_FIELD_VALS));
    rd_cg14=new;
  endfunction : new
endclass : ua_int_id_c14

//////////////////////////////////////////////////////////////////////////////
// Register definition14
//////////////////////////////////////////////////////////////////////////////
// Line14 Number14: 139


class ua_fifo_ctrl_c14 extends uvm_reg;

  rand uvm_reg_field rx_clear14;
  rand uvm_reg_field tx_clear14;
  rand uvm_reg_field rx_fifo_int_trig_level14;

  virtual function void build();
    rx_clear14 = uvm_reg_field::type_id::create("rx_clear14");
    rx_clear14.configure(this, 1, 1, "WO", 0, `UVM_REG_DATA_WIDTH'hC0>>1, 1, 1, 1);
    tx_clear14 = uvm_reg_field::type_id::create("tx_clear14");
    tx_clear14.configure(this, 1, 2, "WO", 0, `UVM_REG_DATA_WIDTH'hC0>>2, 1, 1, 1);
    rx_fifo_int_trig_level14 = uvm_reg_field::type_id::create("rx_fifo_int_trig_level14");
    rx_fifo_int_trig_level14.configure(this, 2, 6, "WO", 0, `UVM_REG_DATA_WIDTH'hC0>>6, 1, 1, 1);
    wr_cg14.set_inst_name($sformatf("%s.wcov14", get_full_name()));
  endfunction

  covergroup wr_cg14;
    option.per_instance=1;
    rx_clear14 : coverpoint rx_clear14.value[0:0];
    tx_clear14 : coverpoint tx_clear14.value[0:0];
    rx_fifo_int_trig_level14 : coverpoint rx_fifo_int_trig_level14.value[1:0];
  endgroup

  virtual function void sample(uvm_reg_data_t  data, byte_en, bit is_read, uvm_reg_map map);
    super.sample(data, byte_en, is_read, map);
    if(!is_read) wr_cg14.sample();
  endfunction

  `uvm_register_cb(ua_fifo_ctrl_c14, uvm_reg_cbs) 
  `uvm_set_super_type(ua_fifo_ctrl_c14, uvm_reg)
  `uvm_object_utils(ua_fifo_ctrl_c14)
  function new(input string name="unnamed14-ua_fifo_ctrl_c14");
    super.new(name, 8, build_coverage(UVM_CVR_FIELD_VALS));
    wr_cg14=new;
  endfunction : new
endclass : ua_fifo_ctrl_c14

//////////////////////////////////////////////////////////////////////////////
// Register definition14
//////////////////////////////////////////////////////////////////////////////
// Line14 Number14: 188


class ua_lcr_c14 extends uvm_reg;

  rand uvm_reg_field char_lngth14;
  rand uvm_reg_field num_stop_bits14;
  rand uvm_reg_field p_en14;
  rand uvm_reg_field parity_even14;
  rand uvm_reg_field parity_sticky14;
  rand uvm_reg_field break_ctrl14;
  rand uvm_reg_field div_latch_access14;

  constraint c_char_lngth14 { char_lngth14.value != 2'b00; }
  constraint c_break_ctrl14 { break_ctrl14.value == 1'b0; }
  virtual function void build();
    char_lngth14 = uvm_reg_field::type_id::create("char_lngth14");
    char_lngth14.configure(this, 2, 0, "RW", 0, `UVM_REG_DATA_WIDTH'h03>>0, 1, 1, 1);
    num_stop_bits14 = uvm_reg_field::type_id::create("num_stop_bits14");
    num_stop_bits14.configure(this, 1, 2, "RW", 0, `UVM_REG_DATA_WIDTH'h03>>2, 1, 1, 1);
    p_en14 = uvm_reg_field::type_id::create("p_en14");
    p_en14.configure(this, 1, 3, "RW", 0, `UVM_REG_DATA_WIDTH'h03>>3, 1, 1, 1);
    parity_even14 = uvm_reg_field::type_id::create("parity_even14");
    parity_even14.configure(this, 1, 4, "RW", 0, `UVM_REG_DATA_WIDTH'h03>>4, 1, 1, 1);
    parity_sticky14 = uvm_reg_field::type_id::create("parity_sticky14");
    parity_sticky14.configure(this, 1, 5, "RW", 0, `UVM_REG_DATA_WIDTH'h03>>5, 1, 1, 1);
    break_ctrl14 = uvm_reg_field::type_id::create("break_ctrl14");
    break_ctrl14.configure(this, 1, 6, "RW", 0, `UVM_REG_DATA_WIDTH'h03>>6, 1, 1, 1);
    div_latch_access14 = uvm_reg_field::type_id::create("div_latch_access14");
    div_latch_access14.configure(this, 1, 7, "RW", 0, `UVM_REG_DATA_WIDTH'h03>>7, 1, 1, 1);
    wr_cg14.set_inst_name($sformatf("%s.wcov14", get_full_name()));
    rd_cg14.set_inst_name($sformatf("%s.rcov14", get_full_name()));
  endfunction

  covergroup wr_cg14;
    option.per_instance=1;
    char_lngth14 : coverpoint char_lngth14.value[1:0];
    num_stop_bits14 : coverpoint num_stop_bits14.value[0:0];
    p_en14 : coverpoint p_en14.value[0:0];
    parity_even14 : coverpoint parity_even14.value[0:0];
    parity_sticky14 : coverpoint parity_sticky14.value[0:0];
    break_ctrl14 : coverpoint break_ctrl14.value[0:0];
    div_latch_access14 : coverpoint div_latch_access14.value[0:0];
  endgroup
  covergroup rd_cg14;
    option.per_instance=1;
    char_lngth14 : coverpoint char_lngth14.value[1:0];
    num_stop_bits14 : coverpoint num_stop_bits14.value[0:0];
    p_en14 : coverpoint p_en14.value[0:0];
    parity_even14 : coverpoint parity_even14.value[0:0];
    parity_sticky14 : coverpoint parity_sticky14.value[0:0];
    break_ctrl14 : coverpoint break_ctrl14.value[0:0];
    div_latch_access14 : coverpoint div_latch_access14.value[0:0];
  endgroup

  virtual function void sample(uvm_reg_data_t  data, byte_en, bit is_read, uvm_reg_map map);
    super.sample(data, byte_en, is_read, map);
    if(!is_read) wr_cg14.sample();
    if(is_read) rd_cg14.sample();
  endfunction

  `uvm_register_cb(ua_lcr_c14, uvm_reg_cbs) 
  `uvm_set_super_type(ua_lcr_c14, uvm_reg)
  `uvm_object_utils(ua_lcr_c14)
  function new(input string name="unnamed14-ua_lcr_c14");
    super.new(name, 8, build_coverage(UVM_CVR_FIELD_VALS));
    wr_cg14=new;
    rd_cg14=new;
  endfunction : new
endclass : ua_lcr_c14

//////////////////////////////////////////////////////////////////////////////
// Register definition14
//////////////////////////////////////////////////////////////////////////////
// Line14 Number14: 25


class ua_ier_c14 extends uvm_reg;

  rand uvm_reg_field rx_data14;
  rand uvm_reg_field tx_data14;
  rand uvm_reg_field rx_line_sts14;
  rand uvm_reg_field mdm_sts14;

  virtual function void build();
    rx_data14 = uvm_reg_field::type_id::create("rx_data14");
    rx_data14.configure(this, 1, 0, "RW", 0, `UVM_REG_DATA_WIDTH'h00>>0, 1, 1, 1);
    tx_data14 = uvm_reg_field::type_id::create("tx_data14");
    tx_data14.configure(this, 1, 1, "RW", 0, `UVM_REG_DATA_WIDTH'h00>>1, 1, 1, 1);
    rx_line_sts14 = uvm_reg_field::type_id::create("rx_line_sts14");
    rx_line_sts14.configure(this, 1, 2, "RW", 0, `UVM_REG_DATA_WIDTH'h00>>2, 1, 1, 1);
    mdm_sts14 = uvm_reg_field::type_id::create("mdm_sts14");
    mdm_sts14.configure(this, 1, 3, "RW", 0, `UVM_REG_DATA_WIDTH'h00>>3, 1, 1, 1);
    wr_cg14.set_inst_name($sformatf("%s.wcov14", get_full_name()));
    rd_cg14.set_inst_name($sformatf("%s.rcov14", get_full_name()));
  endfunction

  covergroup wr_cg14;
    option.per_instance=1;
    rx_data14 : coverpoint rx_data14.value[0:0];
    tx_data14 : coverpoint tx_data14.value[0:0];
    rx_line_sts14 : coverpoint rx_line_sts14.value[0:0];
    mdm_sts14 : coverpoint mdm_sts14.value[0:0];
  endgroup
  covergroup rd_cg14;
    option.per_instance=1;
    rx_data14 : coverpoint rx_data14.value[0:0];
    tx_data14 : coverpoint tx_data14.value[0:0];
    rx_line_sts14 : coverpoint rx_line_sts14.value[0:0];
    mdm_sts14 : coverpoint mdm_sts14.value[0:0];
  endgroup

  virtual function void sample(uvm_reg_data_t  data, byte_en, bit is_read, uvm_reg_map map);
    super.sample(data, byte_en, is_read, map);
    if(!is_read) wr_cg14.sample();
    if(is_read) rd_cg14.sample();
  endfunction

  `uvm_register_cb(ua_ier_c14, uvm_reg_cbs) 
  `uvm_set_super_type(ua_ier_c14, uvm_reg)
  `uvm_object_utils(ua_ier_c14)
  function new(input string name="unnamed14-ua_ier_c14");
    super.new(name, 8, build_coverage(UVM_CVR_FIELD_VALS));
    wr_cg14=new;
    rd_cg14=new;
  endfunction : new
endclass : ua_ier_c14

class uart_ctrl_rf_c14 extends uvm_reg_block;

  rand ua_div_latch0_c14 ua_div_latch014;
  rand ua_div_latch1_c14 ua_div_latch114;
  rand ua_int_id_c14 ua_int_id14;
  rand ua_fifo_ctrl_c14 ua_fifo_ctrl14;
  rand ua_lcr_c14 ua_lcr14;
  rand ua_ier_c14 ua_ier14;

  virtual function void build();

    // Now14 create all registers

    ua_div_latch014 = ua_div_latch0_c14::type_id::create("ua_div_latch014", , get_full_name());
    ua_div_latch114 = ua_div_latch1_c14::type_id::create("ua_div_latch114", , get_full_name());
    ua_int_id14 = ua_int_id_c14::type_id::create("ua_int_id14", , get_full_name());
    ua_fifo_ctrl14 = ua_fifo_ctrl_c14::type_id::create("ua_fifo_ctrl14", , get_full_name());
    ua_lcr14 = ua_lcr_c14::type_id::create("ua_lcr14", , get_full_name());
    ua_ier14 = ua_ier_c14::type_id::create("ua_ier14", , get_full_name());

    // Now14 build the registers. Set parent and hdl_paths

    ua_div_latch014.configure(this, null, "dl14[7:0]");
    ua_div_latch014.build();
    ua_div_latch114.configure(this, null, "dl14[15;8]");
    ua_div_latch114.build();
    ua_int_id14.configure(this, null, "iir14");
    ua_int_id14.build();
    ua_fifo_ctrl14.configure(this, null, "fcr14");
    ua_fifo_ctrl14.build();
    ua_lcr14.configure(this, null, "lcr14");
    ua_lcr14.build();
    ua_ier14.configure(this, null, "ier14");
    ua_ier14.build();
    // Now14 define address mappings14
    default_map = create_map("default_map", 0, 1, UVM_LITTLE_ENDIAN);
    default_map.add_reg(ua_div_latch014, `UVM_REG_ADDR_WIDTH'h0, "RW");
    default_map.add_reg(ua_div_latch114, `UVM_REG_ADDR_WIDTH'h1, "RW");
    default_map.add_reg(ua_int_id14, `UVM_REG_ADDR_WIDTH'h2, "RO");
    default_map.add_reg(ua_fifo_ctrl14, `UVM_REG_ADDR_WIDTH'h2, "WO");
    default_map.add_reg(ua_lcr14, `UVM_REG_ADDR_WIDTH'h3, "RW");
    default_map.add_reg(ua_ier14, `UVM_REG_ADDR_WIDTH'h8, "RW");
  endfunction

  `uvm_object_utils(uart_ctrl_rf_c14)
  function new(input string name="unnamed14-uart_ctrl_rf14");
    super.new(name, UVM_NO_COVERAGE);
  endfunction : new

endclass : uart_ctrl_rf_c14

//////////////////////////////////////////////////////////////////////////////
// Address_map14 definition14
//////////////////////////////////////////////////////////////////////////////
class uart_ctrl_reg_model_c14 extends uvm_reg_block;

  rand uart_ctrl_rf_c14 uart_ctrl_rf14;

  function void build();
    // Now14 define address mappings14
    default_map = create_map("default_map", 0, 1, UVM_LITTLE_ENDIAN);
    uart_ctrl_rf14 = uart_ctrl_rf_c14::type_id::create("uart_ctrl_rf14", , get_full_name());
    uart_ctrl_rf14.configure(this, "regs");
    uart_ctrl_rf14.build();
    uart_ctrl_rf14.lock_model();
    default_map.add_submap(uart_ctrl_rf14.default_map, `UVM_REG_ADDR_WIDTH'h0);
    set_hdl_path_root("uart_ctrl_top14.uart_dut14");
    this.lock_model();
    default_map.set_check_on_read();
  endfunction
  `uvm_object_utils(uart_ctrl_reg_model_c14)
  function new(input string name="unnamed14-uart_ctrl_reg_model_c14");
    super.new(name, UVM_NO_COVERAGE);
  endfunction
endclass : uart_ctrl_reg_model_c14

`endif // UART_CTRL_REGS_SV14
