`ifndef AHB_DEFINES7
    `define AHB_DEFINES7

    `ifndef AHB_DATA_WIDTH7
        `define AHB_DATA_WIDTH7 32 // AHB7 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH7
        `define AHB_ADDR_WIDTH7 32 // AHB7 address bus max width
    `endif
`endif
