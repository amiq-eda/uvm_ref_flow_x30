`ifndef AHB_DEFINES10
    `define AHB_DEFINES10

    `ifndef AHB_DATA_WIDTH10
        `define AHB_DATA_WIDTH10 32 // AHB10 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH10
        `define AHB_ADDR_WIDTH10 32 // AHB10 address bus max width
    `endif
`endif
