/*-------------------------------------------------------------------------
File1 name   : spi_config1.sv
Title1       : SPI1 environment1 configuration file
Project1     : UVM SystemVerilog1 Cluster1 Level1 Verification1
Created1     :
Description1 :
Notes1       :  
----------------------------------------------------------------------*/
//   Copyright1 1999-2010 Cadence1 Design1 Systems1, Inc1.
//   All Rights1 Reserved1 Worldwide1
//
//   Licensed1 under the Apache1 License1, Version1 2.0 (the
//   "License1"); you may not use this file except1 in
//   compliance1 with the License1.  You may obtain1 a copy of
//   the License1 at
//
//       http1://www1.apache1.org1/licenses1/LICENSE1-2.0
//
//   Unless1 required1 by applicable1 law1 or agreed1 to in
//   writing, software1 distributed1 under the License1 is
//   distributed1 on an "AS1 IS1" BASIS1, WITHOUT1 WARRANTIES1 OR1
//   CONDITIONS1 OF1 ANY1 KIND1, either1 express1 or implied1.  See
//   the License1 for the specific1 language1 governing1
//   permissions1 and limitations1 under the License1.
//----------------------------------------------------------------------


`ifndef SPI_CFG_SVH1
`define SPI_CFG_SVH1

class spi_config1 extends uvm_object;

  function new (string name = "");
    super.new(name);
  endfunction

  uvm_active_passive_enum  active_passive1 = UVM_ACTIVE;

  `uvm_object_utils_begin(spi_config1)
    `uvm_field_enum(uvm_active_passive_enum, active_passive1, UVM_ALL_ON)
   `uvm_object_utils_end

endclass

`endif

