`ifndef AHB_DEFINES20
    `define AHB_DEFINES20

    `ifndef AHB_DATA_WIDTH20
        `define AHB_DATA_WIDTH20 32 // AHB20 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH20
        `define AHB_ADDR_WIDTH20 32 // AHB20 address bus max width
    `endif
`endif
