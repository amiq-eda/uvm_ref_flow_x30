`ifndef AHB_DEFINES21
    `define AHB_DEFINES21

    `ifndef AHB_DATA_WIDTH21
        `define AHB_DATA_WIDTH21 32 // AHB21 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH21
        `define AHB_ADDR_WIDTH21 32 // AHB21 address bus max width
    `endif
`endif
