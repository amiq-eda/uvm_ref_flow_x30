`ifndef AHB_DEFINES19
    `define AHB_DEFINES19

    `ifndef AHB_DATA_WIDTH19
        `define AHB_DATA_WIDTH19 32 // AHB19 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH19
        `define AHB_ADDR_WIDTH19 32 // AHB19 address bus max width
    `endif
`endif
