/*-------------------------------------------------------------------------
File1 name   : apb_subsystem_pkg1.sv
Title1       : Module1 UVC1 Files1
Project1     : APB1 Subsystem1 Level1
Created1     :
Description1 : 
Notes1       : 
----------------------------------------------------------------------*/
//   Copyright1 1999-2010 Cadence1 Design1 Systems1, Inc1.
//   All Rights1 Reserved1 Worldwide1
//
//   Licensed1 under the Apache1 License1, Version1 2.0 (the
//   "License1"); you may not use this file except1 in
//   compliance1 with the License1.  You may obtain1 a copy of
//   the License1 at
//
//       http1://www1.apache1.org1/licenses1/LICENSE1-2.0
//
//   Unless1 required1 by applicable1 law1 or agreed1 to in
//   writing, software1 distributed1 under the License1 is
//   distributed1 on an "AS1 IS1" BASIS1, WITHOUT1 WARRANTIES1 OR1
//   CONDITIONS1 OF1 ANY1 KIND1, either1 express1 or implied1.  See
//   the License1 for the specific1 language1 governing1
//   permissions1 and limitations1 under the License1.
//----------------------------------------------------------------------


`ifndef APB_SUBSYSTEM_PKG_SV1
`define APB_SUBSYSTEM_PKG_SV1

package apb_subsystem_pkg1;

import uvm_pkg::*;
`include "uvm_macros.svh"

import ahb_pkg1::*;
import apb_pkg1::*;
import uart_pkg1::*;
import spi_pkg1::*;
import gpio_pkg1::*;
import uart_ctrl_pkg1::*;

`include "apb_subsystem_config1.sv"
//`include "reg_to_ahb_adapter1.sv"
`include "apb_subsystem_scoreboard1.sv"
`include "apb_subsystem_monitor1.sv"
`include "apb_subsystem_env1.sv"

endpackage : apb_subsystem_pkg1

`endif //APB_SUBSYSTEM_PKG_SV1
