`ifndef AHB_DEFINES12
    `define AHB_DEFINES12

    `ifndef AHB_DATA_WIDTH12
        `define AHB_DATA_WIDTH12 32 // AHB12 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH12
        `define AHB_ADDR_WIDTH12 32 // AHB12 address bus max width
    `endif
`endif
