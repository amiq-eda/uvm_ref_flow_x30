`ifndef AHB_DEFINES13
    `define AHB_DEFINES13

    `ifndef AHB_DATA_WIDTH13
        `define AHB_DATA_WIDTH13 32 // AHB13 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH13
        `define AHB_ADDR_WIDTH13 32 // AHB13 address bus max width
    `endif
`endif
