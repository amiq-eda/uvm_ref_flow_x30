`ifndef AHB_DEFINES26
    `define AHB_DEFINES26

    `ifndef AHB_DATA_WIDTH26
        `define AHB_DATA_WIDTH26 32 // AHB26 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH26
        `define AHB_ADDR_WIDTH26 32 // AHB26 address bus max width
    `endif
`endif
