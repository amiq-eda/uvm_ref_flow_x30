/*-------------------------------------------------------------------------
File20 name   : test_lib20.sv
Title20       : Library20 of tests
Project20     :
Created20     :
Description20 : Library20 of tests for the APB20-UART20 Environment20
Notes20       : Includes20 all the test files. Whenever20 a new test case file is 
            : created the file has to be included20 here20
----------------------------------------------------------------------*/
//   Copyright20 1999-2010 Cadence20 Design20 Systems20, Inc20.
//   All Rights20 Reserved20 Worldwide20
//
//   Licensed20 under the Apache20 License20, Version20 2.0 (the
//   "License20"); you may not use this file except20 in
//   compliance20 with the License20.  You may obtain20 a copy of
//   the License20 at
//
//       http20://www20.apache20.org20/licenses20/LICENSE20-2.0
//
//   Unless20 required20 by applicable20 law20 or agreed20 to in
//   writing, software20 distributed20 under the License20 is
//   distributed20 on an "AS20 IS20" BASIS20, WITHOUT20 WARRANTIES20 OR20
//   CONDITIONS20 OF20 ANY20 KIND20, either20 express20 or implied20.  See
//   the License20 for the specific20 language20 governing20
//   permissions20 and limitations20 under the License20.
//----------------------------------------------------------------------

`include "apb_uart_simple_test20.sv"
`include "apb_spi_simple_test20.sv"
`include "apb_gpio_simple_test20.sv"
`include "apb_subsystem_test20.sv"
`include "apb_subsystem_lp_test20.sv"
`include "lp_shutdown_urt120.sv"
