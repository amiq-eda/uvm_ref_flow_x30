/*-------------------------------------------------------------------------
File15 name   : test_lib15.sv
Title15       : Library15 of tests
Project15     :
Created15     :
Description15 : Library15 of tests for the APB15-UART15 Environment15
Notes15       : Includes15 all the test files. Whenever15 a new test case file is 
            : created the file has to be included15 here15
----------------------------------------------------------------------*/
//   Copyright15 1999-2010 Cadence15 Design15 Systems15, Inc15.
//   All Rights15 Reserved15 Worldwide15
//
//   Licensed15 under the Apache15 License15, Version15 2.0 (the
//   "License15"); you may not use this file except15 in
//   compliance15 with the License15.  You may obtain15 a copy of
//   the License15 at
//
//       http15://www15.apache15.org15/licenses15/LICENSE15-2.0
//
//   Unless15 required15 by applicable15 law15 or agreed15 to in
//   writing, software15 distributed15 under the License15 is
//   distributed15 on an "AS15 IS15" BASIS15, WITHOUT15 WARRANTIES15 OR15
//   CONDITIONS15 OF15 ANY15 KIND15, either15 express15 or implied15.  See
//   the License15 for the specific15 language15 governing15
//   permissions15 and limitations15 under the License15.
//----------------------------------------------------------------------

`include "apb_uart_simple_test15.sv"
`include "apb_spi_simple_test15.sv"
`include "apb_gpio_simple_test15.sv"
`include "apb_subsystem_test15.sv"
`include "apb_subsystem_lp_test15.sv"
`include "lp_shutdown_urt115.sv"
