/*-------------------------------------------------------------------------
File26 name   : spi_defines26.svh
Title26       : APB26 - SPI26 defines26
Project26     :
Created26     :
Description26 : defines26 for the APB26-SPI26 Environment26
Notes26       : 
----------------------------------------------------------------------*/
//   Copyright26 1999-2010 Cadence26 Design26 Systems26, Inc26.
//   All Rights26 Reserved26 Worldwide26
//
//   Licensed26 under the Apache26 License26, Version26 2.0 (the
//   "License26"); you may not use this file except26 in
//   compliance26 with the License26.  You may obtain26 a copy of
//   the License26 at
//
//       http26://www26.apache26.org26/licenses26/LICENSE26-2.0
//
//   Unless26 required26 by applicable26 law26 or agreed26 to in
//   writing, software26 distributed26 under the License26 is
//   distributed26 on an "AS26 IS26" BASIS26, WITHOUT26 WARRANTIES26 OR26
//   CONDITIONS26 OF26 ANY26 KIND26, either26 express26 or implied26.  See
//   the License26 for the specific26 language26 governing26
//   permissions26 and limitations26 under the License26.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH26
`define APB_SPI_DEFINES_SVH26

`define SPI_RX0_REG26    32'h00
`define SPI_RX1_REG26    32'h04
`define SPI_RX2_REG26    32'h08
`define SPI_RX3_REG26    32'h0C
`define SPI_TX0_REG26    32'h00
`define SPI_TX1_REG26    32'h04
`define SPI_TX2_REG26    32'h08
`define SPI_TX3_REG26    32'h0C
`define SPI_CTRL_REG26   32'h10
`define SPI_DIV_REG26    32'h14
`define SPI_SS_REG26     32'h18

`endif
