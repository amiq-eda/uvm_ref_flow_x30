/*-------------------------------------------------------------------------
File28 name   : spi_defines28.svh
Title28       : APB28 - SPI28 defines28
Project28     :
Created28     :
Description28 : defines28 for the APB28-SPI28 Environment28
Notes28       : 
----------------------------------------------------------------------*/
//   Copyright28 1999-2010 Cadence28 Design28 Systems28, Inc28.
//   All Rights28 Reserved28 Worldwide28
//
//   Licensed28 under the Apache28 License28, Version28 2.0 (the
//   "License28"); you may not use this file except28 in
//   compliance28 with the License28.  You may obtain28 a copy of
//   the License28 at
//
//       http28://www28.apache28.org28/licenses28/LICENSE28-2.0
//
//   Unless28 required28 by applicable28 law28 or agreed28 to in
//   writing, software28 distributed28 under the License28 is
//   distributed28 on an "AS28 IS28" BASIS28, WITHOUT28 WARRANTIES28 OR28
//   CONDITIONS28 OF28 ANY28 KIND28, either28 express28 or implied28.  See
//   the License28 for the specific28 language28 governing28
//   permissions28 and limitations28 under the License28.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH28
`define APB_SPI_DEFINES_SVH28

`define SPI_RX0_REG28    32'h00
`define SPI_RX1_REG28    32'h04
`define SPI_RX2_REG28    32'h08
`define SPI_RX3_REG28    32'h0C
`define SPI_TX0_REG28    32'h00
`define SPI_TX1_REG28    32'h04
`define SPI_TX2_REG28    32'h08
`define SPI_TX3_REG28    32'h0C
`define SPI_CTRL_REG28   32'h10
`define SPI_DIV_REG28    32'h14
`define SPI_SS_REG28     32'h18

`endif
