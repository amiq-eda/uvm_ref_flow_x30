/*-------------------------------------------------------------------------
File29 name   : test_lib29.sv
Title29       : Library29 of tests
Project29     :
Created29     :
Description29 : Library29 of tests for the APB29-UART29 Environment29
Notes29       : Includes29 all the test files. Whenever29 a new test case file is 
            : created the file has to be included29 here29
----------------------------------------------------------------------*/
//   Copyright29 1999-2010 Cadence29 Design29 Systems29, Inc29.
//   All Rights29 Reserved29 Worldwide29
//
//   Licensed29 under the Apache29 License29, Version29 2.0 (the
//   "License29"); you may not use this file except29 in
//   compliance29 with the License29.  You may obtain29 a copy of
//   the License29 at
//
//       http29://www29.apache29.org29/licenses29/LICENSE29-2.0
//
//   Unless29 required29 by applicable29 law29 or agreed29 to in
//   writing, software29 distributed29 under the License29 is
//   distributed29 on an "AS29 IS29" BASIS29, WITHOUT29 WARRANTIES29 OR29
//   CONDITIONS29 OF29 ANY29 KIND29, either29 express29 or implied29.  See
//   the License29 for the specific29 language29 governing29
//   permissions29 and limitations29 under the License29.
//----------------------------------------------------------------------

`include "apb_uart_simple_test29.sv"
`include "apb_spi_simple_test29.sv"
`include "apb_gpio_simple_test29.sv"
`include "apb_subsystem_test29.sv"
`include "apb_subsystem_lp_test29.sv"
`include "lp_shutdown_urt129.sv"
