/*-------------------------------------------------------------------------
File18 name   : spi_defines18.svh
Title18       : APB18 - SPI18 defines18
Project18     :
Created18     :
Description18 : defines18 for the APB18-SPI18 Environment18
Notes18       : 
----------------------------------------------------------------------*/
//   Copyright18 1999-2010 Cadence18 Design18 Systems18, Inc18.
//   All Rights18 Reserved18 Worldwide18
//
//   Licensed18 under the Apache18 License18, Version18 2.0 (the
//   "License18"); you may not use this file except18 in
//   compliance18 with the License18.  You may obtain18 a copy of
//   the License18 at
//
//       http18://www18.apache18.org18/licenses18/LICENSE18-2.0
//
//   Unless18 required18 by applicable18 law18 or agreed18 to in
//   writing, software18 distributed18 under the License18 is
//   distributed18 on an "AS18 IS18" BASIS18, WITHOUT18 WARRANTIES18 OR18
//   CONDITIONS18 OF18 ANY18 KIND18, either18 express18 or implied18.  See
//   the License18 for the specific18 language18 governing18
//   permissions18 and limitations18 under the License18.
//----------------------------------------------------------------------

`ifndef APB_SPI_DEFINES_SVH18
`define APB_SPI_DEFINES_SVH18

`define SPI_RX0_REG18    32'h00
`define SPI_RX1_REG18    32'h04
`define SPI_RX2_REG18    32'h08
`define SPI_RX3_REG18    32'h0C
`define SPI_TX0_REG18    32'h00
`define SPI_TX1_REG18    32'h04
`define SPI_TX2_REG18    32'h08
`define SPI_TX3_REG18    32'h0C
`define SPI_CTRL_REG18   32'h10
`define SPI_DIV_REG18    32'h14
`define SPI_SS_REG18     32'h18

`endif
