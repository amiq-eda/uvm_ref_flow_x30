`ifndef AHB_DEFINES27
    `define AHB_DEFINES27

    `ifndef AHB_DATA_WIDTH27
        `define AHB_DATA_WIDTH27 32 // AHB27 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH27
        `define AHB_ADDR_WIDTH27 32 // AHB27 address bus max width
    `endif
`endif
