`ifndef AHB_DEFINES18
    `define AHB_DEFINES18

    `ifndef AHB_DATA_WIDTH18
        `define AHB_DATA_WIDTH18 32 // AHB18 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH18
        `define AHB_ADDR_WIDTH18 32 // AHB18 address bus max width
    `endif
`endif
