// IVB15 checksum15: 2692815514
/*-----------------------------------------------------------------
File15 name     : ahb_master_sequencer15.sv
Created15       : Wed15 May15 19 15:42:20 2010
Description15   : This15 file declares15 the sequencer the master15.
Notes15         : 
-----------------------------------------------------------------*/
//   Copyright15 1999-2010 Cadence15 Design15 Systems15, Inc15.
//   All Rights15 Reserved15 Worldwide15
//
//   Licensed15 under the Apache15 License15, Version15 2.0 (the
//   "License15"); you may not use this file except15 in
//   compliance15 with the License15.  You may obtain15 a copy of
//   the License15 at
//
//       http15://www15.apache15.org15/licenses15/LICENSE15-2.0
//
//   Unless15 required15 by applicable15 law15 or agreed15 to in
//   writing, software15 distributed15 under the License15 is
//   distributed15 on an "AS15 IS15" BASIS15, WITHOUT15 WARRANTIES15 OR15
//   CONDITIONS15 OF15 ANY15 KIND15, either15 express15 or implied15.  See
//   the License15 for the specific15 language15 governing15
//   permissions15 and limitations15 under the License15.
//----------------------------------------------------------------------


`ifndef AHB_MASTER_SEQUENCER_SV15
`define AHB_MASTER_SEQUENCER_SV15

//------------------------------------------------------------------------------
//
// CLASS15: ahb_master_sequencer15
//
//------------------------------------------------------------------------------

class ahb_master_sequencer15 extends uvm_sequencer #(ahb_transfer15);

  // The virtual interface is used to drive15 and view15 HDL signals15.
  // This15 OPTIONAL15 connection is only needed if the sequencer needs15
  // access to the interface directly15.
  // If15 you remove it - you will need to modify the agent15 as well15
  virtual interface ahb_if15 vif15;

  `uvm_component_utils(ahb_master_sequencer15)

  // Constructor15 - required15 syntax15 for UVM automation15 and utilities15
  function new (string name, uvm_component parent);
    super.new(name, parent);
  endfunction : new

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
  endfunction : build_phase

endclass : ahb_master_sequencer15

`endif // AHB_MASTER_SEQUENCER_SV15

