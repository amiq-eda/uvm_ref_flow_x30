/*-------------------------------------------------------------------------
File21 name   : test_lib21.sv
Title21       : Library21 of tests
Project21     :
Created21     :
Description21 : Library21 of tests for the APB21-UART21 Environment21
Notes21       : Includes21 all the test files. Whenever21 a new test case file is 
            : created the file has to be included21 here21
----------------------------------------------------------------------*/
//   Copyright21 1999-2010 Cadence21 Design21 Systems21, Inc21.
//   All Rights21 Reserved21 Worldwide21
//
//   Licensed21 under the Apache21 License21, Version21 2.0 (the
//   "License21"); you may not use this file except21 in
//   compliance21 with the License21.  You may obtain21 a copy of
//   the License21 at
//
//       http21://www21.apache21.org21/licenses21/LICENSE21-2.0
//
//   Unless21 required21 by applicable21 law21 or agreed21 to in
//   writing, software21 distributed21 under the License21 is
//   distributed21 on an "AS21 IS21" BASIS21, WITHOUT21 WARRANTIES21 OR21
//   CONDITIONS21 OF21 ANY21 KIND21, either21 express21 or implied21.  See
//   the License21 for the specific21 language21 governing21
//   permissions21 and limitations21 under the License21.
//----------------------------------------------------------------------

`include "apb_uart_simple_test21.sv"
`include "apb_spi_simple_test21.sv"
`include "apb_gpio_simple_test21.sv"
`include "apb_subsystem_test21.sv"
`include "apb_subsystem_lp_test21.sv"
`include "lp_shutdown_urt121.sv"
