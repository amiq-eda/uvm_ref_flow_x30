/*-------------------------------------------------------------------------
File14 name   : test_lib14.sv
Title14       : Library14 of tests
Project14     :
Created14     :
Description14 : Library14 of tests for the APB14-UART14 Environment14
Notes14       : Includes14 all the test files. Whenever14 a new test case file is 
            : created the file has to be included14 here14
----------------------------------------------------------------------*/
//   Copyright14 1999-2010 Cadence14 Design14 Systems14, Inc14.
//   All Rights14 Reserved14 Worldwide14
//
//   Licensed14 under the Apache14 License14, Version14 2.0 (the
//   "License14"); you may not use this file except14 in
//   compliance14 with the License14.  You may obtain14 a copy of
//   the License14 at
//
//       http14://www14.apache14.org14/licenses14/LICENSE14-2.0
//
//   Unless14 required14 by applicable14 law14 or agreed14 to in
//   writing, software14 distributed14 under the License14 is
//   distributed14 on an "AS14 IS14" BASIS14, WITHOUT14 WARRANTIES14 OR14
//   CONDITIONS14 OF14 ANY14 KIND14, either14 express14 or implied14.  See
//   the License14 for the specific14 language14 governing14
//   permissions14 and limitations14 under the License14.
//----------------------------------------------------------------------

`include "apb_uart_simple_test14.sv"
`include "apb_spi_simple_test14.sv"
`include "apb_gpio_simple_test14.sv"
`include "apb_subsystem_test14.sv"
`include "apb_subsystem_lp_test14.sv"
`include "lp_shutdown_urt114.sv"
