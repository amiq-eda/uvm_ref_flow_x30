/*-------------------------------------------------------------------------
File25 name   : uart_ctrl_pkg25.svh
Title25       : Module25 UVC25 Files25
Project25     : UART25 Block Level25
Created25     :
Description25 : 
Notes25       : 
----------------------------------------------------------------------*/
//   Copyright25 1999-2010 Cadence25 Design25 Systems25, Inc25.
//   All Rights25 Reserved25 Worldwide25
//
//   Licensed25 under the Apache25 License25, Version25 2.0 (the
//   "License25"); you may not use this file except25 in
//   compliance25 with the License25.  You may obtain25 a copy of
//   the License25 at
//
//       http25://www25.apache25.org25/licenses25/LICENSE25-2.0
//
//   Unless25 required25 by applicable25 law25 or agreed25 to in
//   writing, software25 distributed25 under the License25 is
//   distributed25 on an "AS25 IS25" BASIS25, WITHOUT25 WARRANTIES25 OR25
//   CONDITIONS25 OF25 ANY25 KIND25, either25 express25 or implied25.  See
//   the License25 for the specific25 language25 governing25
//   permissions25 and limitations25 under the License25.
//----------------------------------------------------------------------


`ifndef UART_CRTL_PKG_SV25
`define UART_CRTL_PKG_SV25

package uart_ctrl_pkg25;

import uvm_pkg::*;
`include "uvm_macros.svh"

import apb_pkg25::*;
import uart_pkg25::*;

`include "uart_ctrl_config25.sv"
`include "uart_ctrl_reg_model25.sv"
//`include "reg_to_apb_adapter25.sv"
`include "uart_ctrl_scoreboard25.sv"
`include "coverage25/uart_ctrl_cover25.sv"
`include "uart_ctrl_monitor25.sv"
`include "uart_ctrl_reg_sequencer25.sv"
`include "uart_ctrl_virtual_sequencer25.sv"
`include "uart_ctrl_env25.sv"

endpackage : uart_ctrl_pkg25

`endif //UART_CTRL_PKG_SV25
