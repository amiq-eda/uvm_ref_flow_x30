/*-------------------------------------------------------------------------
File16 name   : test_lib16.sv
Title16       : Library16 of tests
Project16     :
Created16     :
Description16 : Library16 of tests for the APB16-UART16 Environment16
Notes16       : Includes16 all the test files. Whenever16 a new test case file is 
            : created the file has to be included16 here16
----------------------------------------------------------------------*/
//   Copyright16 1999-2010 Cadence16 Design16 Systems16, Inc16.
//   All Rights16 Reserved16 Worldwide16
//
//   Licensed16 under the Apache16 License16, Version16 2.0 (the
//   "License16"); you may not use this file except16 in
//   compliance16 with the License16.  You may obtain16 a copy of
//   the License16 at
//
//       http16://www16.apache16.org16/licenses16/LICENSE16-2.0
//
//   Unless16 required16 by applicable16 law16 or agreed16 to in
//   writing, software16 distributed16 under the License16 is
//   distributed16 on an "AS16 IS16" BASIS16, WITHOUT16 WARRANTIES16 OR16
//   CONDITIONS16 OF16 ANY16 KIND16, either16 express16 or implied16.  See
//   the License16 for the specific16 language16 governing16
//   permissions16 and limitations16 under the License16.
//----------------------------------------------------------------------

`include "apb_uart_simple_test16.sv"
`include "apb_spi_simple_test16.sv"
`include "apb_gpio_simple_test16.sv"
`include "apb_subsystem_test16.sv"
`include "apb_subsystem_lp_test16.sv"
`include "lp_shutdown_urt116.sv"
