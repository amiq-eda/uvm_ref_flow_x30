`ifndef AHB_DEFINES11
    `define AHB_DEFINES11

    `ifndef AHB_DATA_WIDTH11
        `define AHB_DATA_WIDTH11 32 // AHB11 data bus max width
    `endif

    `ifndef AHB_ADDR_WIDTH11
        `define AHB_ADDR_WIDTH11 32 // AHB11 address bus max width
    `endif
`endif
